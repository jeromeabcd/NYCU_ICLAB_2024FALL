`ifdef RTL
    `define CYCLE_TIME 20
`endif
`ifdef GATE
    `define CYCLE_TIME 20
`endif

module PATTERN(
    // Output signals
    clk,
	rst_n,
	in_valid,
    in_data, 
	in_mode,
    // Input signals
    out_valid, 
	out_data
);


`protected
H;,#-BNLH&S_\].A;2)ebfUD,01J./2+9</I-C/[Q)H;K.;9X;:d,)5K&@>J+=<7
#@T]O7)SM]6#G<<&#<P_I<[TZ^LWJgG]fI)6e4S.]WKA@2P9;6&M7+6+8.35N<Q4
/FR?>\T3eHBZ?)g-J=,2_BIcd)^C;O+AJ9S<<M^T9bdHYA9?2A/ZZB8@(Xg9::Z\
S=CDC#7GXMdd3.[XYFLB_SIc5$
`endprotected
output reg clk, rst_n, in_valid;
output reg [8:0] in_mode;
output reg [14:0] in_data;

input out_valid;
input [206:0] out_data;


`protected
@aR(QBFeEB(P0]6W)O86G(JNX8SfHVR2<9)GdZ=Z]&V&].&=ZCG;7)GUY9.d5H-G
f>:Y.HT,;>OSXe,eX.Pa(1-ALYK#1R#RRA7H:11[Z)Q&28g@<bFBR46N9G0deN__
-eQ2K=3>P2;_<;<:7KMLKQI42/Vd##6b;^BIbe:7FR,[8+9V@TC@=+<N,c[/SX>>
NHLS=:dJ1VVGObVB]5;J-)683HMYPR]2<?(\B(99=1O_c<0];Pe>?<0>Y=XSSV\]
9B4;?]254BCMO>FXND=Y(F,-f,35=0cS[g+Y&AZ5b60eXTC^1bSS>Fd,deYLaPaK
LMg>?<<P9:KHZ+;HB0aYZQ/+2P#KM>YK,3>=0_10?77J<&>gJIWM&gZVUMHBeD/\
WeJ#I2af.:,gUJ8e^\^U0&.>IS,[,SO#5>cP]Ga-@JO-HN2>?H<<\J=9C][?,5,K
]ZOFBUEf,Q?K8b&]/47AF5QV_.[gX\S#6R>PA(a/WKLL[9[dM>,<2^O?Q:6Bba@@
b,TbL2Dd[=G0BJR__>T-/IbY]g#W.,5</+HI-HJ8P[W&FR:A?45ET3)bCeP#.HBg
-@K9cGI^?b(2eO\/,]da(Xg2YNYN,=Bd)\_VZ&&NK8db1K1DQ]@deK)=X@)>&T19
9H0?c_e@?8GU:4,FF)3521f\C->S-?NFP3SIL7VCg63GT/PJY[25V@eL<I/dT[bR
5\:SCea-&3Yg8Y[(Z@L=cQ&EU3AFO&E(_B;HH9(&TM;230\>L-?/U[5TJG&?Hd0:
T1d3c&8/#BeV;(<4C-IbGR>DPI^QFKN1I&B.[=[&[-D_Y&MM=>]Q:Y#fQOV4dTH6
88+fNg](f>ZaBBg,eNKE:UZa)WZI?67OB0:B#U^HT###.Z^^bab0<R8]^1CAU5#J
#G]H>\DcN@SS@LgI1XED=T2JD0g+<S2IBYSEZdCRRKM3HYQQXXfCZ[eVWcT4MG9L
Ga2Sa4UdB1dRJ4]>gK:60]AeDB>M82FG0QV=NK/8?O>C_XPG-\JN(R6>?++0@gd0
DLS+GCH[&63U3?6eL<GY>GI;K:P3&DE^DA6QP.abUN<c)=+IdTNQ\JWLXM(\>XM>
d2=?Dg>.8JDC4VAE+URWI8e7)V:M3BM]JNY@^AFbB0F9XY#I^c[>XHQ5LL/6A.fQ
ST\;05(,@XI)(<&-\M\MEc>faVV37N7Pe]W()0#=]]b2H+12(M?1Ib75>TW8VB@G
;P2OgN4M1RU3-.IaWZ4a_FGe6:??bMddg=O@<&E4\?N>;44eT)^-_b[e:a=gJKGM
SVcM0[g#2e(^?B>;B-PC&\[[93US?LCK#DC>:<9ON9@0HSX1D6@\8CTHS.OQ63EK
0]gH6SXFG8TbLO##<9M_c\5ebDg-L5&@5(eL+-feN?^GP1c182&S=#SIfgbY0<+^
(;_/4d4/H5(^8=+b/HIdER>/+Xg7d/g4ZgSJ\DB^#<K5;7[@1B9,E66O#/,A7P^-
dG0L^-2YadVN[ITHUP_4VF7\dM6#+XE&KK[>KbS/\BMb0TbI<H?UR+:\Ye6XVELE
GN[I76/M3FV4QRC[2]^_S4IA@a/ATCdK]\eQDce8ZgfN_XSG2d<eX+a,A_D&0&P+
ZD4H,gX&>N[6WY-N)Z(EOa3I_gX8&(8LJ1b73\bg,,<g&4:4Afe@5_>1T_<N<be[
YLOB?1TaCSVU+e-7#.G86MRL-NHEPO1d,GcC;9CDVdX/b_RT49\b[,.e5P.FC@6-
^))\79AS829NRF]HKgIR=6[&(7UKSZU4e<26aS(+-UHaBf8TY.0ae+I>2dgBO>RD
39(FY-ZT()N-]I@&bHPLZ0:17V+Z;G1Va\F.GRNU+K0UK)CX-Y;g23DMddO73D()
U&Qf5L?4gPJ>8B4>(f=[?33:MBAI2WK9#>L&5&Y:ceTPEb0e0=<>Y6CZ[HL(d\3P
-;LId@:16;;;W+F=ZY&aC.#6@P-<(#dd:g@+L:bQe9SB.@^=X2D8;SAbC6.M81XR
?]Zce1&(e3>63/P5V7P=f?T-,/MB_DPI6RDGH&XU79;IHOD]fVUH6(F)C^#Z3feZ
\.fEd8cfH#7Te0+_8[FMSO@2O/>X0_3^:U,f66fRV@-ZMF_&XeT>daLa]-c/de:@
;SC_&S,FP9FK1b@Z05V]B7?5b\EUa_bTJW>V3RH.+cE:Y/[eJ22)F[RfC=Tc-fHG
c+XBe<1TR:@^25ceY#(4TL#HX>OQEL6aPH;FK#OH#J]5T>=[dc?22&5V&8(MAOHV
FW)@/<Ec7=BO9CFR+#eN-eN0.-+,R#DE7D_1NUL_e<QVXXE14/C[7J2(?CDV)_>d
JC;3:dD?_I)&BVNE,^Bd9M6ce)_+e9dNN\^dZb;Y6:26SA?cA2a91@RJF/0XRE:T
^2X=C&QMW<bIHF2SGWF>4LCJb>E25&+@&,_&[JZ0FV1K1C2Sb0g+-N-M)AH1ZR.;
CO8&Zgc-TE1c&ST2AX[VE9.fI0>77CNcb3CfQ)QPdEN?a+1A/2VX)65YO:LXLdE;
.>J+Ma/8VY]Za@?=>[-(XVCdZB@K\3<AE&HO,L<P3FRVOB-<S;7)3UTHF+H&W6P]
-,N]Tfa-PY>0TaV4e>LdJ4YLWGa/A.MN.bFZ-;2DSYH//NG+6+7A/cT4Be):L#P3
CDJ,D<A?U=??.#7?7.bNP8?;0K+1,g2H</U5J-J/d]5e73V+\D;&.Q.WL(AfP=EW
1(MV:W1I#M7S+_E(\+</9I[(B[/\+X6OCFAC^aVSP:<+FS+eBKDSb/)S0c=+]DW1
Z,dT=V)UGS@3R&TR=_Y4VecRPTgB_8#S4U=<H7eR?<QOV2F.9>[+[_AdSVPJ3XFK
[E(_>3F1B#J;[G4:/WO?79)ZQ/2)GfCbGH>_YYR5d]Eda#D6Z./I4Q_]-JN7P(C;
FJZ&cAYFYa;Ig<6fg^<J]bGR(Rf#.A(WS-aaRE8P6P5MZ_4Wb^J[O3X>UWNd]YWS
^eeOZ6M[SBDf2fDI:L#AY[;caT7e-HCJ>TMLadTK+Yg/UVGU1Ra0fF\5;G6HR#(B
JG_,H5-MU4RQf;a1WRbOD<-)?DT2PFS;R>T\JBRIMdD/>VFC&C:0@<>&C@<\W08b
#RY=Xg2(YKSAKBF/W/_BOM-/Ob]UX98cN4b#3-+6eZg-Df:X6SKR8\S-bU:f@=N:
9ZF2USWY14_.9C\?-We]TC?)D>329W24V13&#,Dg<XS5X?N2#+SYL1)1c870>6UB
#GA._[,TPRSS^aBN>?X@F)KS<;XbXZD^SCG^O+-+-AbE_FM_08V05X5C)K&H5//L
O&cA=HbLd58]?aS_BVUQDV1gSfNO0PDUKI;d=L-P4KPg6X;K:1QfA>NP\KI:^8J>
B1Wb&bQYJG^@U&>#>bfC,>[BVb=__;@E27E:b#\\<WSA0MbQa&7WP&[:PbRFLce\
\Hf>C6_WS(]baNDGdcP?I1?=>MI@()H=&gOb9>2W=ab_8)SJ()/HG7P#\/C;+PAb
BIHY(@0S4)_7d<.6L#M83D;\H(_JY(\0275c6/G\GMF[R-G&K#C#^F<:5^T0?8/R
SaEQV9S)0E+R#H[X0,SNK.X?BHEP&F^Ye(OZC7KUd.LY/81+4(;,@&.7/A.QdfMF
Y9-EV:;)CbTJP[?13))N(]5C&c/]0RWdRbZA@F&7J.:0VMI0KO#;4[)^M+H;A6H>
+A1&eE5c+LN^GdH]T0Df>\5^6eO/A-]27+TXNW0Ndf[;FI^-14Ma&ZA<8H/XZ<Rd
]#&1H^:K@eE9(VGP1C&OM;>@/&VS,H9&8:&O(8+PV7LBVA/4#)AgMAgL>W-/Bg55
X/Ga65OQ0H)CD,;dDK4@ZLZeGHPZ26Q)AeZ7_0D-^WLKN([D8##]-;6JM;/E[/8.
_[B(V.(6ES\Mb[XgS91cFU/:-?CQG\LO.gW.#gX;PT-]HGM1\,[e\a61AKZC#^^&
.]\([S/DC_:P@)HPZd3(7(^d(B:<2T+IgU_S9:]\3<N/-M<)KWA9dZZ11eKLRZ(@
)c)_:[.S.I04O6<@dAPKG@\6&NVD-MXD0bQFYRb]GIK@.SXgN)A\KZ7<K_8WWgR1
fK19(IPAYgd:)Y)>B.@KH;P?Z,P;2+gP\e\)\Y57WVJW^,:Ya=X\XY\:HQ73MB<9
?)=B>2g^03YZe,#Fd;BT8B7>C;EE5[8^L4fR0H2T955X]2[VeaY^24#+P)P8T5^/
#?R@Q85c._I8@bYC2M1#6-)/[?;fAKXU=(=:QA(LS<HDH@6,1?+6.SP3OFJ;da3@
_Xd8L-&&E+eO4D#8A.2HDFgA@dI]>5.[cF;TS:(]@ORfX3&gBJ);[L3Wa6MN+L]a
PDU>cFcUK\OV+YT,BP@dLb>ITNaXRaY#c34^HD5/@/4U-;HO7A>85K9+O-W,3M##
@-dTKUXVHA_=C45-Z9eX9N3B]=TC#g9L)EGX[gNfXI4f0c@90AZHV.[71(@686)&
0ET6IOGJ7OG..-T(/=ZYSAR9GQaPe;#8HG6f^EMJ07/Ue81\]A-+J\da;R?5b21b
\eLgdb3E/b>DJ+S92YULbS7g?]eb\J4#EQ8Z-/\E#VA,1FH2(KR[\e+T_)g?X8(T
_31C[@a>7R=N,MALW8L@/9K=AX9]V(77a+6eWM2?YK9+FHDV:9:]TET>1U>f<LOS
;6AE;C<=>M;aC3RD7Oa+>2Q(CV0GA[G>J75LA<+d,ZS\<\H:;#C>4GZ@aVICV+/(
,8NVgf]M)E^@?\?76-4G(06=>@cZOC-R9\?+<Q(NBCC0T;/FMfU9HRJQGISAO4^F
N]:dL8ac[9XY>J:Z?G49/YFELCZ73]NQ8T@aNWd6YO0/8(C.cTZ@/3(A04J5_)R&
+EB/-R1@_73Gg&NP>R8BcH#E#N+SeMD#7#:6&WDP&XeUE]TdQ_^BB9WA@C9_P?X;
e<AM?\c#QVC,@;ZO5LaV+>/LWY+1RH@PddR+O-I9?@9AT<1R7V>S<ER0G\cgDP(E
c]A#P\Q\#b-6Z5;L.@3E.RDdP3A\2Od8]QW7S;#,Vd4>DSZ2Y;8eH]gaNFJ\XdS;
H6/KX09]+Q?fT5W-C>[W/>FEb8[1(?bN,9?ZRS/g#]>C]<O@U3\X&f7NISdf[JfY
FQW9Y18f7P,Y5db:f8c<g]Y[SFg#(+Z\X+PFdd0>55.a>/<O;4Q-7BcS;MH#D7-)
g6)27[MV.aRNeF9C?+AR>VO^H&SM83LE5@I^A7e1=EG&+-L7dOZf?E1J05D4<^S9
0(?=Q]4=[&ccdA[EBBR=NWG-eOATIbKQEES@5:(KWM.2Yd9;f)]Q)Z8Z=,)g;Q@+
D<5K;,TD#MCGJa\FDcQ3Nc[Sb[0Tg^EM-aK4]KQ+bMI8W\M1@eD8:Z86D]AHIJg;
3FNX5DG=M:M-E:f4_\Q(HU92/];EYJdRc8R\==Q[Y&,\W+>81QJd4Zb]9d\VO26W
B0agICg3XdE,3\#B4@0@)(WA(N([1\dC)P3E3F_QET@HU]A8d>I>NLT>C+HacS,5
QfKB/T-^;(?aUa,De#-1bDg3=Z2?94A9/H-D8)[?EN+6#:,4Y+A^c>>V0+U<K6dM
+g,H1;-g8(c)02[+NdJ2Z=fZd\e4RdVVL-;E)#&C,>>8^GFabVRAP/P:cJb.ee]d
=P4H?I/NJDD4<fE&a2:U?3G?H4X9b4=[0V=VXg?VHda-&EKS1C+&(N^\V2c53;^P
QYg=gJ^,&N;bE+V<a/EGfaT9E]d3[6,HR7-M[bI+Jd&6cFb;B,]bY=I)Q@K2QGdc
P/cNbf^OVM19WaE).\Kc&FGGVGggCc-[.#@d[?RD4Z-T6@C&.AdA>9\<Rc&UY?QN
(@7P:R0BKW<]_4a?-J57R9d@UXD/<A6AZT:YU(+Z(&@(We.d526D,GT6^O9+f];L
R4/.CR3?=->-T]RNP@5085.B5b8fF@?7T;eeX]/]S/W&2NcY,[5/DSf&0fW9D]1\
8_Z:NBMZf1(FIENENO)/X[F4#I2YA,P9,7MK6;e7?BYB)AX1d#fARM_OH:SRHVA]
V).cI]I[6g)@FAP;L5^OYf1P?^6X8F[=<<bEL9+Mdb&4DGNcd<EYRS1;@dX3Yf@G
e\1aL@+X7a94-91QaU=-MZZ_W8-Oa(d3eY9;W7GI^THU,T+.)fB^d)QJGbYSB@gf
Y].cP(YEaKgZe/H^\_Tf5;A&43+dJC?7K2fPNQaW^O3^=:?ZOb]Oe8#Cd0>)TQ8X
\76K;?0dFK,+e;@65_0KHP15(8DOEZTf_f^g<eSeW;HK:3dfODR82I^33G86Pbc9
d6:IKVJ(DQA>Z:O[6_<X)EU<=P(&_>8#dcE-7?(2cbf9?aY]TBL_O<>,&D29V4WY
T7I0[/[G@[TeSH_MI/ZgHc0#F^<PdZ>[AF1R4ZcHXR/(6T)?JdJ42gd56Y(ZU_HG
00]>/,1Q0C^R&56]]&g(8SZGGT/-:J&A+OA+APeQ>3L06Y>6K/<X>ca\IAe9MU#c
.FT]40HS3L2L=OHR)M3:=:&&P-a>=3gT@F,A;[Z9-L3e/25MW/W8dDg3Fg,OW@)C
dY&(>(,;&VL,4L<]-KZH8f^-VgaQ&T8^YIG#Y9b>IOa)2G42DK7)Q<:/#ZAP\9NM
Y\/:#P.FIXP8RA;8UT(>La[Ef#g6V91:VTb_6QTJH)3P4IFN(GdgP&6Y6&6/,F8b
1E0(b9gCPORK/fVD+YU;JFYS5X/fEc-(-^/=612/8FVF77@/PR#TYP13Bf>GN-_>
W0O\7.e?.[HG03/dE#O9VN\:CX6^C17+2,68V#b5Y^SY,\6A&)aZ7CQT^W(X?d->
X1BEDO?R/f5#6SOQ&DPU2P;eQ>H)6#FO@U?AIaMWc4Y3O77^[=(B:1ED-BMQW3.6
F7F^A-32)T;72-(TY[gT&QL;3Y1(UAP.4_L1_cHAW;ZeI.0&<W35GJY187#X.P4g
KF6/f-8OP/]2bMGS)afc#J76B7[L=(/0;UYdMJKK?/T&=3:WP)2GY4B(,Uf^2-:>
8EBOaMOIM(NTfYY8A/RRSP+W@B<QH:g+\9T?F9AU/PGJ2=G00Yg+O=4A^cK7afdG
M.^H9Tg?G@@OO>>HGV+##U)A.]CN(T?\gY&Ec>Iaa=SZZ_4SK:Ze[OW8P6CFFMSJ
[.3-87Y,Hc).VH2^:PW?)O3Zg7gQKeMJeU?dM:)9S[^GEdVe,:a8_e/QAaY,H4T-
6LG@c)&68A67CP9dB#3cHG5>)AO=H7XMAb&ADBBPPF&YK&UUN<Z.U2)[0Z#cH/&P
D[[HD5#,3RgANId/&b+_G#FS(GG:P1[d^ZEbe6b?FD4,12D4SU)a:;ELW7@b?6,4
K:J(/609aE\>#Z-FdF5LHLc?Yb@2HcN8B7SRX.Ra?##KGcUHLYEI@NS]/[GK1dXZ
^)e:eEU#2eW>LJOd:LXa.8CYOVU_R5A:?JeI7;,3<DV\5)bPcVbCYKLQ/ICGMGNJ
GG^H2FD4Q&HJ]#M<T[Vb?V9EIPD3N/?[dIaOJ+R4IA:PDPWXS2R8)90+R>aFWfJf
IbNLV]Q][EG-1^P0I=#N7eF&dI#K:?fP>-TcbRO2c+TH>F7<60P#B/e(12LLe#IZ
5.<=^N+#NWW5&)eH;.1L?;D+IIWS4Z#.608[72OfJ-T_1CEF&8U<Q=&VFfL/f1^>
3<0)O],]O]JC&XeYN.)W#eS4@L,M<MgC(-]R<Q+2ZOb7g,@LQ]AQS+:.PPe,SNJI
>.H3Q2X5b#43H,05L8TA2HF(]NPW_Q0g@LXYXC/O[gX,GA]6Z5G_[aQ1VaK@=6_7
d1<BK0f1:YF__;K1(L:8@5C;aF9-2JQcR9B9[6Q1U=VX)J^VDg1/OdUAF\A@=TQN
<bg;<?a]8UM#?(1IA>]SUUTA>EM8^LHRg2JV7DELR1g)=9B98OI0R>,3XFa[RL1a
dCDg,FZ3KMgZ/aO:>,ZPZD=<N\KH\^?-Aea_S(e?9D2Ycc_d97[d6[DYTPWCNV(4
-AO5][9^,/?:CZ(5R.4A_=48TKfXRXX[e4d&\NU;QE(6TCLV8EPO:?T)KRQgTD7I
_9H:EX\JI8RX<].:Na6:F1gE)/.(dH+JQX.CDMbd:9&6.7F-E&2,SX.Rd+0.B5bW
=F+DR>/163_4WWeG3H0/=E8KRJ4XH(KM1g>,D4RgZfb3.g+83_>8/Waaf.4MecU;
-MaE&0EXF0^H&V]e(<1&.?eH4TV<,:f=daY2O5Ab:IC2.gN15T#.OK7Zb4=2-KgH
[W8<AEX<A>2Y)3@4UC5ed(<4d<aQbLMKJWJK<?<C5d]egBb?8KcS6a^,<+fE^?1X
b_\P6\V2OaH@Nd]ZME^P(+[TeM5U@AE#M@VVQUQdAf8[S#+B?O4]):1=H_XQR4\X
\#a.1GZU;5[^WRD<]3@;7&.K_:(6M<:HLcL5[_?a5Ne7.BKf_E+A,Z7PJ9A=2U;E
f/]\JQ-0HM7?D8-459Y:)Lf^@=T?D(4?>9N^OX^5#e6QZ=F)PQS&K9K<[9gQS.Z5
g[10)58=UL#-C3[7f1<ZLN?+^HfB+ZHaE+H^@e([e(+U&5&82Gd9@R1.XVC]MJW?
Q8(;HJ6^Ce\T15J9e&#)PD@Rb<ADJI?^VNWA15)H4fJg4>>J+D7T7]Y+(3<NR,6U
;OCHPDU_NT64A)Q,Z)c#^DE9DG<>M>@P+B)8).RM0HJA&=UT&GagX+5^;/P^7XKV
3N=:)EQIWUBJ8XSOCfT=>RD_?KDDE#EPVP5GBD60@Na[X@d)c55Z=^Q5)&RFA9W1
C?RHCI0Od253Y+C+N11Ub@/TQ(N++CeC33,5SV3&d1>+c@bdXT:2e?cM4RYB,T9R
<DB#W<,Dd8bg+\3J7=P1eIKeRIJg&L>//3>=Z51UE#B+Z?8Y]733F6#_.I/[fX(\
-(XK9UcMB.,LGb0&_J).F5EEHAdIcfa_>P^)RP->1&b87)-fMPLL\&cXRHca]&2b
5R+a^Y-O8X\8&c1aVX2VRa2]JD)BGW\6ZHOJE-MD22bM\>Kcd5RPOLdHS^:N7[cU
15J0=S57PZHT-/Ee1MWI5;,eH7d#&ZZ#<W=3TRb\)3=R&K.ITJ?+S^)#,)M.+0:b
(@b@-HW-@>ZA@A89\\H\M(Tb)M;I8UQL@<f4=9@1NO)#CN7BSL6Pb-07Fe_&M(ZA
JI<KQ88_SZ#RN8_(I-[]4S:K(9]^=_TO+A&@=g7#.C)]3V1PJQM]1=&ABG[8+c:f
O=;.PPbU8#KH4S+A^CXBKd5,P3,<HLC60MaCF\WKJRW(G&QIGf@TDd_0Yc:0eUKI
GaYYPLb,J]P#^#P;;FDP8&#5I3/aeE/)S./1MFdF^3(>UMIWTV<Y-J0aLVIJ,YK^
XX3B4M6EUWEbJ?AZHbTf6\H2O@B&O]Q3)#KV:->V]:7_Ga]Kc,)>4YGNEANg1NRS
g^@a3@5c9^JCW7WXeK?=8O7NA249_I4S44G]M=L:cPI+a2X,QBGcGG3^#1-LOM6)
.W_[LQP0R]g32VbHPIfc?Tc0#_J&PNeWAA=#/RRY:1&[:=X/PPfXZ&e(<?M8KZUF
c(I2KeQeY1Q@J^3<QJFT2cKG\CL7)<B464Ha#:a]Z[+8@c<]T4WLE2?_\e0_>,Z\
\NQF::Sf^YdUdVJ7=W&;RN5DA#F)XVR3Ka?O7</[GZOU+;1DJD2L3EN&MZ=2IUeg
JXa6AD\]#QQ/PGEDCeN2W2(S;-a2]YCBc)1J7.Mg1=W2O_AfQ5/FO7#0PTW(=MY7
ASQ=FV.c=K+gIV2UUV;=E#,?NK/?cO[V0bfg<;\T,FUfA<@O[4/gMWR/O+VQf1#J
IWU84,2P6XJc0OQZ1)00OU7\1Kb#X?c#dWH/=PW?1CQRg743>/EYDOCV\1VT)4LH
&,,PRT^B8UOR<He\\/9WbL_bU;#Jcc,Td_cgI7,^_NM,?3+(W]4Q3D.3+ff,E:/X
2\K/W.ZN4HS89@?Ge.](::1S1.G-;/]\YF^N9,U3\dcWHRTL<7C=6EL3[XVIMBgQ
)X=T5,WQ&9P^XQ,_+[_3VBd393I]eAT5.8^_S8KJZLVGEV>L2T<CEb56L>BYG-&Y
BfffGLeCEJ>LQKRTP+8,OM/UEdbC4OL/@bR9a(-dG83c\MDcGdbKV.K?OMQ4@[?Y
,c;VXN6?T=,D]&R./?OB(:V1JBAXZ?E(6BJ81CZ.;Kb@OF0c5]XF=\UY_D62eR?U
+3A(05I:b#=g<cG7d8DW(+O[@e[dQ5<g)W8=Ma0H7+1=4a&YNDc#FCeOba&^S,,S
gFQG8I5L59R@\5+_Acg:8;_6AMbDL],@-T]fBVSgF1,YTBJ4C(O_bH<T-bgP7N:B
>7XE+]>53_T5DLRb#HXV;.SXPN(B5<S6^QWY2P:cH4[N0@\e;5)8BQIB1]c.7>]N
)d[L&WTgc?MZYB\_2P+JecR_W>f/HbEd6>W])=S<Lc=#g0_-eBCVVG)?A4Yc&,_X
^&J>J4d8[eP\WZ=&O3U])aD8-.?AQ^ZI1ga5+8V&gAJV\ZbI<(BQA5&JF-3I&\2R
R<VeO=G]gK@>Jg8]3]D9-OAC;0F>HG_b#JDO1K1+5g97#egZ&Z4:?ae2WPX6eY3-
A5bM,_H5T\HBL>\S6=^g-SX8=C/8)05QK;]B=ZPE<UJ.3I]230P:U<(PQ[NL88D<
,^GV4/>[WT[F4RU/OaWKcMeMT8D=^T4S=;JgS2NA8\1)aVS@RMD&fS;@J]HO)eWK
UGF<g;XGM4YI/Ec^PUaG]/V^(^5=AXNe/_I/X3#gGCCW8/\YDb[M-5T+#2GK9,Ke
)M<7eY.JP)F8]BeWHbE.YRgBO78>B^JZ-83cY^ZLBTB>]HZ1g3f4fgN=A:-1/1gB
&bE;4\a_\U28YV]A5b79FAG:c#?W_Gd/LM30G#M?<:+&f7=.&^R&PU(ccdH_<FT.
)^>2JI5BJ-b2ePY>dKY=DCW)=+/T:&(O>_OgdgSK14X;35@YAXOSEdJAQd1dY#O\
.;+6fHcbB\W;]8Be_H#:fb#bK_VQ/c?]d5ZL[0e3/F.O:0aWJXMLLg]XJ#?.R+,U
7L45B3EWK8,3EG:HN,cP&M<]=A;Q+HR=>d/N8fIDP\H/f6S0+8H<PHD:.8W8I47;
8N7X^eVR/]#S7X;D(5C]0LMJNCe+/J=6>(:(]+0O-K>Y.);XNXA&_L&TV>>;G=@I
&[0FZCg9:&2^#.9@Y<?R5Qf+@9W50c1@O3Fb8.KCUGH.D@()/Kc])MX?bABe[-4.
&U=SCfL;6->Gf+Ba1G<TX.3^0C/6.aV5fZ3VMD_4LOJ#527+UP=YCPM^@W[f@BWd
^&N60aR+VgSY6#R:Q&+Ia&25G;fN>R_&N86;A06@Lg^^dIWOG6+;J\=KN)&ce.Hf
ZH6a7[J3&g/EdX99\&SYX1K5K-<[Ac]62a5.Nd-<^FY]_CE3O^:1:.X2H<aZ?ICB
VX4f_&5GgDD^?KG)e1OB;TfM,Y)@/fTH>C(B,1(\&b-gX8>XG^N,TYH^690c+c3#
IF]De)VX]+QAeZeB/0Q,IPB5aJ7.9X52RZ9Kc1&,#3EQ-(+82A1YKbF=>,9NL4CY
(^=G+<S<[OaT7;DP61BVbEC,)S^8TG_b[>&?A6LB-P?CHWN64dW\O/A[(BTU&JNU
Wg#Z4\9N2eb7;_(U(#?RDJU4eZDCRD;#QI3&fcOK[RXB,95FHf7Z5U1@X?T[97cW
L4JH#/NZ0N^2<Q_P,1c/@+V<4PC8YZAUN\d:&E.LRO_:BL+5G-aTFW9eg)gW21;c
^GdIFN70A(W,dN8?F;\;GZQ6DRR0K4de>TSA&fMAg#CK3FW/C5[,+71D)@?b@3CO
LT[]G)RN8<,;^@V-A,6,g=QTWUcMICIXUIIQFA9/5S<O/P(Ia>eA;:^9A_]MY\M9
L:H@P=+-A8?MFJRcWD^/3f6]gTGZ.f7P7;?aTdA,K>?Q10WIN?>V_]APQ?0ad<U(
,_Z-L_A:3M[IU,a9\XP.1&/@fM2I>X5;a,3Q6=Z=H>McZ+W;@_U<EBRFA.dBP/]V
99IU=]Y-F0;.Af;dMgA5P76^#GN[&HVEDRK[[@;B<3,P&E(NF[:HE/(;QJdCe).?
T/@)Oe-UU#:NE;45ABA2F9WPB//a,J_QM)#V+X,N/CPP8,_=X06EJ#?JGJJcIN.4
H)01?dDb82P5N)IY:P]-]P=6bVNQ(&I6T(.bILA)aXgZQZA:^^WM90R&0P6]IU[5
&O/E1KS3cCVYOHOf22P-M4g3=]#:PPMR?&S&S8)P1\;c7(IRCG8K5I,\JFH\30=9
eB/ED+6)/2MJY<fRZE]>e]?Ya&=E]HZL+#D?-&]PK/_^RH&Y,=N#7-;96)Y00)[6
\R6#^UI=3f9ZP&c7G+G]1(0[7(S+?N_P0UYT#[fKa4?(Q]E+NNZagK>O4c-,SbK]
7?TbWGUOK:-g\Z(aa)^P0bD#>EU+Aa:2>9AC9C)e\c3#I/#9&HC<<IgKLB2X(:f_
6ILe4FS\A,/I05-<N)Y-R--NQC8Sc>U_CQIR:;ZV_\4G_eecD>07^RbCY+aOA#A/
8a6<#RJY=YfK.C4PI]@TT<6.-&,4.Z22L1?BGAE2N6LZIEG+-DV<bIbUOGK&^.D>
Se(G.Kb4:4C6KYGA]/9Cc]M22J3^cTY@OB_<Y/^F)]Q16)==>E;WA\RC1b>?DAff
&:5TEgGP7@_YC#B\U5H(6)OTabY.-A,@1+6/D8d7f)e)[BPGRHW1?0H]c]K7LAET
?;U#bBOAYM8/FNQA3=U0:JM\+EA+be:bad):@(VU4F24a@K#]K/e;GSPa+0><3L>
=e]:#R<f_0Q(fL9V2Z8:g&.gF(a:,,_B,ccBCR#J<Q^Q4W/6?KG)d[O=G@P]GYM5
4GD\OLfN)IW7=23LMRE?-J@Z#@)R8_N?/G>[(K_RYaPT[Y:^Cd=@]SM4A+.<8^(U
+)JS:]_;&]8/:/\J:XgEH1K&fF;IS]=BY^OAK-_./c);3TD@cN^EcZ:Y+(^7<GAY
V.BAaU#7&#-)Y1#LW@EMG79I+7JJ8./eB=>NF3KZWeX08;Z.Q5M815[P^])=g^AH
==T;a8HSRI0_P#]HT2FI^EV@R3IAM;)_O^/X#,-:N[;@<Z:GR&Y(eO.29W::f9:;
OQD+NTUESZdC:Ec9IQ\XURgeAS54?)e?.dJQe58?LX6caAGQEE:Ld.gZ>.]^2Q84
2gUBH0bb-^]Da7Gc(OVD:M5KE-M&X02F&8&[:PcM2SO.<EFYT4<IXT(YW1WC&B#_
B)FID\=YJVV=4D1[_5MQPcD]^2]c:CG[BPKFQC?L0b\8JgI<^-7C3Kb60:1Q/HR2
2g,,J(M^B:@8@E9ZB[Q<DKaI^A>:dSQI.2Me6;MYF3(;Mb5VI@B;Z_[Z=e8<9?fT
F3B,Gb(P8^2ES,K-K>?H6(;U,:H;-WI8)?+\-)b82O3@0AP&b[g]V_)E)?@/36XO
>C=_^gAb1fA9bRGR(Efe8ggK#J]>dQZ_SEEaTH(^(8#9QUfW,>E^c.2M,L9NCG)0
6CaagW=\.\6<+;bR>@aC:C>+LU#<X5WZ@;U+6K@,-6FJgYKN+T36IQQdeG^a>A2f
>-@,#LL&Tc.GX]#Ac:gce]L8>;BVJGd>OWVfbRNF5A4cK.I@>?=:81#<2[B#TJI>
VcU\@[(EFLe18F_^[a_.e+S@/&9]A>H/CWW3a2BBPd=1J^Fc2Zca9WTOAYc056PP
aZ-EF;];_+WD.6ZX(W<LSX[cYDaI(BaaRG>[XJXBQFEC5BO#WAU<QNIG3PdUCZ.#
5G7R_\Xa5XP0@JcFgJKe:=2Y.#=Zg)P,6SES:e.TGYTU^0]#+e;@T\(g.N)?dS?S
4G]9^&4P2/e+2e;Y),3#@CZeLAS>Kga,;P=+/MK&5R8Pc@4#C;[:MI6gKZI;1OJI
=^<.DDUX3L1bMFOU)WF</F5NPXW4Q)gSH1bHW8FePg[74QPQ<Y6ICVKUG]/JO2QQ
9g5Y3b?>7NZ5Y^Ldb1a7/eL2&(\H)[3>)2\[(^Kg9QTID>N:;D<06CY;J(@5H&X/
XXPgR5]_..S45W?+M.-)(FIF9aG\>>/GNg.+@GS&M=?+[^;Z#K[KNSUI=-XM0R+V
D5;]dbGWKS69PELG)86IYUCe8A/Xe<2f906;KE]@5,1LA)&H4[PP72+^3QR\e5LQ
<O;<+:X]TS0OaQfb6DcV??SBNNA(R1[4A4N7gQ:<f(GN,;a4]D_^)SV<:Vc0bUR3
4G[:8JMdR4\&C[6-Cc^T<dEJ<IIDQ,7TB:TRT\U@eN:XH&BdE-3S@7ZL<E:3N#>9
(\,6Y_+D:&>9^eaHCXD56>WLcG3?\@VYa&@6d=905AP.Z>]+V@W_FT.WJ3^W=?3]
[V/__-ad9Le4d\<Nd)dNMW:DW4<-3\&XL-]FD196:7ZEU=?ZAC0eg7#)/<EI_e82
5K8KW;McLJ=Ig./2c.FYMJ@H/LD^Va#d0.>_LE<\^8Fg7J6R.M8MPR-(52fA-gJ1
]Q:=eXF,X&K-8>876cSf_GY]-;:#(G+14[_KJ//4I^Gcb_NOSRPgg\G6f@8_\I&F
4e.)J1#baZUH#N/b+Z6g])fX76S97=W(BbZLf\I9Y+SWD6[C^Y.\&T)@/WRMZ>\5
Y?(==UR7L47-dI^R=5+LWPL)N;-g7?#MdJ0aTOCC/]GUbAB<M]=e//7/GK_BN,Zc
9JT=&]7K,.FXf)-9bMO541]9a0HJGBQ\VZM@/@4OB7gVW3HXe^GIVZG)[=0G8OGS
-=);Jc[J0S,[R5+VC@<8E_,gLRfIWaA8RLW7\-UMd=D=a<CN[O(>6Pe+,,JJcR?/
THb;b9bEN<3>Ve6MDP0-5I,72K0c]<JUeE)f)JMG?Ya)E-J&R1<3]1@aK91/L3dI
001(D]GTNEa,&f+:2GH0_b3=OMH7b&\RV86IANcGQ:)[g7I8[RKWSTOL@eTPD/[;
?6b4[[:+A.:DeD>#.Mc4@T<H#,<SV7cC-QdDXI@+FWI2<S_,6_<1V[O:OQe62^6G
gNE+U_1SQOLVPSbb<#A>B>Ya2-HP3<e3_IPe1#:dIE\?8S>G_M\O0\VcT;+T,N/W
+gZ-M@DRCY<Mf?,UEeFg?P&:8ARL,^\?SCM7O/:DcaJ)H#2:)2MGAB^1>;3a50VT
0e0I/+gF?QUbN<dKAD3?8RNJSWDH1OF>Tb=17NSD]9)Q-[P/W=??OcMNB._VNg,0
?U(9gX0_.5gWJ=(]S,B-ag_/9#25M6<:])eUP_6a-<]bN8eM:EUB[),21=_(McaL
R\<UW2;D1JZU]b\UBA7L9]B@.9PQDCV;#<3KdMc-5)SLD8^TB+f@_;G_8D?FS@C>
KCJGWZFZRA/T&?&IS@I2fMB=[R-,TVMN5JZ10MSNUIC:V?(Mc+VRe:TUG61]K(4(
H5YR#B+:NbE<=:<#H_[60Oa55gSU)SZf[?;GLNW-O>WD,5M<1-\c<1RPR-4-TbZC
gB1O27EX#_E?;?.#,cfH&0BDQa#.RQ)DXCaC.VO3dP][W\f?A@[Ag&C-:SbS)6T?
A+g:L2N)DA2]9)X+Q_b2<S06N6REQOD;:Z\321\F^O:9cK;aP)f^>.D9R.]IO=gP
<dRF\/CK,:WK];60IW<K49>J=R-AVKF/;C@)=ZH=JS=6\&8QKTe3)<^(eD#@Cg6H
HaGFS9@FD\XJAbM#DVR&/+CgY9M8NOZWfcXR7g;8UEf)^C&BN(8)-#9,ZE@X.P4P
Rg2?J9)1#Y&U.:]P6B@eZ7=<B514>c,Ka-64B37>1JIeFUKYg<1;I3c\H-9BJ5\W
?WGO2);VMPc<X4S<b1W4F>SbfGA:C=WL+U9FfERVU+ed.98XOD3+U\d4.YTe0#c4
RSe+\.9=\;+;>98Tc.VN=)1#.#34/Vd;GT-W7ZOO;].:=PTTA.)^QG3(<\(=PPE_
^-;R#K)YS/+F4b955>G4@DA&<M,Ecd&-Y6CM1:Y-RZ6f_+BAA&YIAd[P]1\M@.2L
I4FfXNBP<27FIAGW-KLb9/BC1N1-_EY:F#+(GF&-bSE::UYHDAFXO@_WYfeZ>Y-1
eYXfP>#=FE2M>8&7ZJZ9NVg#g:W20e>?HI[,_7/?;d-L1Y>f]O\Q)2^#OQK6;+4Q
UEJPZ-\d@5F1K>#0g/d?TRSJfRVaZR/@3@b#]RSP#+TQ6IdHT:W[<9,FcRe0Q)dU
WO&RC/T_1TT<P0e;;2W<6<5a<+WAV4.HWd@Y3[0?5[4)aHdW.1?D;AID02(2fD7G
Kd;:5,@BM]1-M45U318bY1O8;KLSJ26M8QXT=ZKQF1LD<N.D8:AJQ=&WXa[dMO-I
U9Y)1ZI)&M,9NA_f+[-.)_SP@)R;L;6QW/OZ]Ya.Y86,@DM<]J_^203a=b>B07OR
FbQXM]2UHBdHRCN9I7.J=82O\e9QX<e3-bf-((8];V+O<-Z\+CJ-#e&SWZ@AcVeP
Kc8I5[TcO1O@c#5Da;V([MV=HX6^V9J0E]_473\1OFVCe/#_DcL:9>d/XQeI)]7J
XJ#2BR/Z&V[&6WecPe2\9,dZ[9=RAVYf-[KU-^LM@IVf4M]UG0(MBM9=cO==]F6b
dRH;/geG5e)=?OBU=U9YIB>/<7.ZD+RLLJ32Z#\Nbb>IVJ>[+@C3JMfU#aUT4@.7
PcM]YR0F)/3#P3(76_?E_=/Ec=EFA+,DU3<\=-fH.FXW:bP[OWIb&<I=eJ,30O./
@J;7[4X;/STK#7HKZR.2HN>5>#4,F35A>8SEG@[#P#AG1O@8TC+4HQ7]I3E#5>.B
]<JbcH=,+\?TKD)=.6HDZeGSWFQZLV/I(^N4>53I>9Sd:/X-)[#2&[#>Q9b/I0#9
Ye\)7HaS[ZP+gQ^QSae/&S8@dS@W,4VM,]/10c<&R&G\]-38]Z@M2Z.8#M417[<b
bQOafD.?#73:A?dTcG5BE34I0F\3@f4bD5CKdA4BFQH<BAJaDGZW,0@QH:/OE,]-
QHIQ/@BDRgKfAC@FZ^c7_&<=;+fb949/.H;85Z9>FIE_E><F/UHX^=1T7K810WG6
IJ1F<Y[I[1^--N3+>PCVV7O^A@Ba/^f@^@2&(]RF-<JV&aeLKd=]\0J6eNd\+CX7
RR#S.E2D=+TeN+??AY_eO5IE(Z5\&A[#[)NO(K8=C@R7f>K=CY,:D4V03/W<9BHY
CYE^d8E0@8V]0)[/1_Yb/;8Ec\]IMQf0MVWaHe&[SC2@UVL;XLc?_&.A;f:SQEF]
MgKW^?gOKDR6a>Ib46WLQ7B^M)^#]D4]dWG,MdL]A_GFJGe[e^)R9B;1SXQ\@,<\
PF9[&IgU-Y33#CDGdZ<.TK.,<,K]D_c8M];b5>cYYDb@7NO02A#VJ_6c;\G2[N_f
3[?JOP5T\Tg16>\ELBfEJUGL1>]83[S;5.dY:2RII(0aGVWT,IEDJP7AddQ+.DTL
2NJZC/S0^Fg+gE9KDA9D[&56DU:14TCI]G(@+SQ]66b(Wb/0>:L9)0(>WNSZ^&S=
dDAC6_N,+aB<16WY_IeB>X[[aFd1DA(Wa6=D+1M7B<J+0:/RY)#RG\HZ:74_MT2b
E.B6CL\Qe.W:,LSPTa2H>@2#=<0ZCSD)Hcf-d[MdCG>[&dC<7YS-8f4]KcbMH6RW
6L,-=aHM2N4YGE2&]ASTHbP9_PV9D49E-4F+_]G1\[CQJKYN/_#?feD4PQ9a=OIJ
gcK(>Q+V5E_TQ]bd&#eVVP?JSR?QK:A[W<80G^H.H6/P=R_5I/@]#IR\c^<_LSeU
5,0:<D;KZ>)S=QQ8X;E\c,6XRGd70[\5g9+04b-]PAaCH,Q9+LJL?L@9=6gC98J8
>R+d,fCRVCN,1^W#(<[\007TZR=<]?_L<9(+RU4T6VCbg5SF-8F4aDID7ZDJg1K,
M2LTWMR//G#BU@QPYJ.,1e9+RJ(JJ7a6-+<@_BUX1b9=UU/^Xg<37.TIce#J9_=7
LS.Q#3H38+?MJ07Ve+T2d9EH7NO,9b4.aI6L#,S_N@;fAY6KO>Jc344.QF,H#88a
[^HIVL2-Q3),JXES,&eQfY=8550J,GDRD/c>E_=N9Wb2#3F66@^<^\K:()E.54@;
\-,@@.FgH(MYfcKO=-)V>7MP]J<0C?NBPK5GaR2ZcP:feN[4e)VLe1H\0;JTH\;Q
1XfFKJcE/RAb_+2VHZQceP&g;J60Q][[::;B]X;N8RJ]@X-.&OK]S56\fOFIN^fL
,MC89+:b)g96>P.H[I0==/(OSZc5<)9;SZQ6P:U=,&E&c&&C81D=,\GB[;2;,_87
b@ZEJ:\[3e<IHW1?.EXI5SP>61d84L_Dg[bXY(f:@9Z]2A_:XW)g0V/:7EY)Pf<4
7O+3L<\4^EHBB:YCbbIY+@S9BN3QPa)2=1)-:gIU/9/.NMCU@A[I38V7FX40(gNK
Te=2L-?OE-1QI4118JW@8]af8]2B2Q:XfK<Y^>8-g:9#gJ9-f@#DF5bdS\SC7<_b
U:7\DE:._-0SLJ53IbacAN^79I_2;VYe4^f>Z)Te3M=K5B86ac/)Pb9?ST#e^aVK
YQ01HM.N.NW.I8LJ(,0A84KN[RB=Gf/_#YTc18=+-5^4L9aY+(S/SFTAB3g5Qb=S
K-(5A5=g:-d7:TD)>OIK07\3/1\K-ZfcQ5G_]P]bTF,PFYdIUc0aPU7&/8PL4VCR
[81@f\b3SX\9CdJOAW2(D6D+NGD/fcCX)[NY:W9?)72M926L;[@9E>(R>&gXFQJ&
S4M3;^ff)Xf6N5bUH?>LfAP4D(REVA]U582V1V-Qa1ZSNL-(G:G<2Q=SaOXEAEX1
UK26?R5>MI/eEEcUD#I:.b,[/e06d^Y)1LRKG1B?1bI:MJ57D:?1dW2gHX65L31=
ZP/<3F<a&<X>\/.FRd)O-?eF)N\-=?AG:86^A\2ZQe3(V1Uaf)CD(Pc<D.c1O\c7
<#dFEV#4+a=)U-@WNCY1D548UNAMR(0cU)&0_PFJ:UYZGUAK379D+J6ERP@\d&](
8Y..MQ<2b_/fa&\EbFLQC#?C:0SVX9,f1/]HFOVY)S8//:D)EN<@f+\GN_5cMON4
Q=;9Ra?R]<#KH=FDOLGA8)PF:Rc\gM/W7AZ6[6UY6#4g7bM:KKQQLNI<BD(N05Y3
=4b6UT>Ib_3[(<dc4(ZMAW]82/U?@R1e<XV3M9;f_P^F:EgDQ>LM2X<[W+N[b-b2
2aQZ/,cf(6^99;Y4d4Y]?ZYRRW+I(Fe[Af;BEXWcR9:NcSS?b0]c^&1Z#/,MW:>=
Tc],NQ4US>bRT)N.g[#cEA0<X@&JRHQ++PYAdcOdA5dA/NFS_\]2M]a.H;IVU#S)
+WgWbOfNT&J]G;Id^]bSaE:OKIA2&U8YO:J<7ZDF049J;3LJ4De=0X]_?J;UE1-,
W^T_QZ.A^=&c0(2Ug)N5(N396AO>8C8JdSA@>#;TBDZRKFSJE]],g/;)X61-^KL7
0/U>RE?+M(H\_LbOCK-5^9:#@KW>NT1H\CYQNYX:H0\H?@4A(-?WLQW5&.\a0T(:
K,^e2CddQb503K;IX)b/A1dGU[FPZU\_[^c#H\8TUXTH+WPNV-(N7F#d92bcC[1Q
Wb.MG7&?C>HGOBe&^74GGG#?+2/C5@WZQ>)7\_-M#GBX6C8#<@V9<ORKcP<\]:AU
/CO,RJ.]4;#VEJ9;a\K:M[?B;]UJD-(&1R8Y\W,Vc2T.I#U;J.ea&O-ZX2VMX^;A
T]LNfY:;_9S]&):XC<[d(T1:F[<\/R)a&N[3f=/E]L,8,b</ETD5&12F+b1/.->:
1X]1FXWD0<+B-V]A>M>+W@1IIYIA#@Ke900V_N(QK=<Vb,>IFD>5=D+.=f9N5NP[
BdbV-@^ILGRCWc/&VD&I2#\RcN421(NH8D(518#]C2]MXaN_LF(;LQT/M0HaU?OW
Hb,NP)5bWe/#I_KS>2@g)#@,7fT]@_[)aYT)[g>;GbbUe&4BM)0d..U_DM#8]\AU
AO4F[)NQUIBY#//aBEF0280--?[5/T_=CHJE869_e..b4KdfMD7be:05cPeH5Ub1
NF@>L:RG^41@Va#UR+K8GJ^JVE8EC[JSC2<]=d4MbOC+_L>6&;.[>f=OY=:ZKcDH
0^@3KK,37X5WEQ,#S/C/S\,KY7,=#QFVX0:^J>#?eQF6/]/]Y1J3O]3e>F&N9P+e
IdcEOA3I^Qe&^3X&QJ-:;Z8=7a8O_4LSCbCJGOO<?Y4I3eGU=37A=NTB]F_SdB[W
.DTH_J=OWe23PQC<5Yc5]FWU/LD?N,X5CHfW#<&-Eba-FYgF/a3LV]P3CSG6aPQH
_a?7CcDT[J(1@E>5#fT):W+?\a;>U8)TbN:3#X.HA:a;K5Q-DdEA[7]b@e4W+LfZ
I7#G9O&I0^0BU+UYWT6R/@SAT8>->e/T;Eb7J(D26\T+#700bP8DG.2c^1G=]PD^
<:B]FAb.#46?Af/f]\&1^M>&fWf_5gXF[3(<cFA#(XV\(QeR>_/a2X7><&M7A-6E
V0aF@H]Q)[.LbDI.dC/=1Z2ICZ#XFDHd61#bLWgX#].1:D3[K0ZZ)I3VW<?#@_\3
:;_TKJ;YeWS]#PDe\KC92[+J_1::VU^)Q5g5Ha,VL4KcHB^8O-SP_dVL_8/]-8A,
?Q0g+GHbDfKb7L-??#E.&e3d^CAM+2\^c.b<Gd^;/U61M.;CPWH,H6I[,;1?:R=,
ObGgMYVbIW7>Q+<;F>08CC4QYIHDNQ;9XdC-RV1Kb5\\_Ha<X<ZB,1VO;KJ7^M+W
Qe4.HG<(76:M7-](K?3G?17S;A^(;6UKC[Hd/3X:Ub_#:4CA&JRD3VPT6<4dBZ)Q
&5&@6X?N[\?.AScJM34AT^T]c4+BZ\KY^Q-T5V4JYedK>N(_G9E<?K<I91)d;dO=
QPKVXR=J7LC1\JKcc=0f^>OV70aYNb+YSGR-Ac2BI<K\dF-A0,,C@IBR,KS]58P;
GP?2O^C4?5^D9V9dWKPgCbR(2:Ag,a[]G<CS>XbI8LcI_a?gP\?^C7-NWL/K5RA3
-Q@7S.Cfg#@-/MQPg[c2KND90C#f/5U\S?:08.,4@,1P)1<?d,2_HCg+I8eWc#Rf
U.5bH[TdP(D:J32TC2R4CZW/bbdabDD#\1#1ARV<_N/QT(Qfb=;B;WcQ>_Je6>7d
X/^Y_Z_@TVa2;UD(=K)e7M&1EK9TN,eM@;_M=44WARH?VT]@\<X.\1eUbaC,:LT@
>K=HJO2MaY2bY35CQ(-LF1[G.L27S)8#RVIS?P/C\+(?=SO4?0T_K5#MM,2I\3,T
GdQG>e]5@6^Y-PQJB=JF[ObM7D/ac=5VEJ_Ib\aA45?9UL&-UK3>ZH^MFMO0;D6Y
=;Ig\GJ#:[V)R/gKJ2R-4L-KO;V[B3I?Qb7V,+A6@QVN>=I464fb(4(65^3<+1[2
IX#JZ1d@1:#-;-Z[UY&8.EZa\1WQ9&W,]cf3,UgNAC?&a3MW_)D(AU[,RbA[0-FM
+^.;C]BN)B+PQO=YDgQcXB]@9B6J/2<DB@af+C#fY@>G[8&#//N?B\3/+1IK@K@[
81=e-=:<f\cHbOXD6_Ga]<SO2L6?+C^;?MZ0T&F8:5CBW;XZ,BMK#W8+1L:4^9XJ
G:ZVU5-[OYP3Qa_^/,NLUg@/].gJb52G71=_0X&:6-=4L5TfgCMJN>E65K\X3</P
D-OHK&].FBgf^)bDA4650&_J.M[CM5Pa21(#g:P&UC&>V:>Oc5RaX40V1Iae@AD2
[f_N_X#X8.SQVP2/ff>R8HC?]&K^YID9<W,6Y&fME#6aLe:XGgC<D/)[[1b>>M-(
[,94VN-\e1Ed_\,ReZ1bNX7@6a9I(#-K)N8-eXLS-UL2bRCA,ReUQf[]SE#01V#Z
]5R0b+EP2@N]/g<9W),#-LdRZYgS(N5@TL1?YTO;@cJ8Y[LA#@2NTSAOFLV7L5(_
[-ENZg=1HVW90ZI4\Bg:dWIe6DLI\R/^]OB4^VY:YCC8FZe.bVC<a.71F;OX)\]&
U9L3_D34egX,DNPROFVE87JY(#:;1d@4WJU:/ZRIN<JFXC87,#ggP5SL3N=L,b-=
W\d+J5-_XR:0J^L3\&&1=a??^3O2S-:O;JY)834:A\KfAQ=Eg?;YJ)SF7+P6Q:PE
/g&5>?HAJ9fJSH8UXB):9@J\9>+S60D:..;SW[2(/^DQ9LP.9d0G&Q7gOH;JJF9e
Hd2@H]BJE/@Xe85Yb=7-_)FRDUVE^6)6JH+9a0QS^4db855EM6+7YH-N11;WWH#S
E@NA&NL#cf76R.8B0bNM0Cc#Y;/Pdf5d/]]?d6O/G#Xb>U3@d+>)+P3\V@FZ71CS
Ad05/7G_.:C/3,)eC0&16gJE+9eaeH\RVe[\#_.B2W<eJ]U(5HI1gZGDL(a;02\b
6\).#JWO;TUYT4RSR.US\_K++EWbN0R,/-ePSc;,aI]Z9DQBU6([3ff9]+f67]#Z
9H?99-;g-HQK3ZN2C_&ZBH/4JEDeLDb,)eD@CebQ_0#Y&f^O9ADZB+TUd8MO3b3Q
N.gF/A&SEBGBY]<#>>NJ,:XJO-XXX]TK]3bLPZ7R-.(=^;GAKA\654cb9;2^bO+H
Y5&)((F-V1TdCdf]NB^I1#gVCcLDbLF.VZ4DM8\K3Ee1RgC[B1#?CSEY]J<AA6:e
AEKC_32L#:+1@SYX2RNXF^0WK/D(aQ^(\M&A]b7&5[8f95OG4:f;9XT0.JU\HPC1
91#G:g3(8U/M1Qfb):H5aC=\]=_/6EHKbYBL:285<ODEZZC[]VHd^3;F<&PcC?7a
.;>/C+3MJ3.<fHXQY+UZZ;5TNTF&7]J9<5L1&\._(C&1DO6b1W5,167c010#(6:.
HXBSMKI,Q98I..H5OR_cEG;<+-Y)J?f966:<-#W>/O4&VCZg1@7EZ>98K7VVHRF[
.DH=_,&/\bUWN7G^KWF#\-@>&L/3b-[NBPe8X_LXUH@H?P,?.ISN.M6^aYDVKTc=
1f9Q99P/N3&BL1[a0gD[N893@>/R_01SC(RWL(OS4F5L/>((&gP?/PdE(XDP_P2D
A52:c4:#@(_5.59#eB93g:a2c[F,L5#BZ&Rc,,;WWY.7eG5E2]=aQT-#aF&WGF.8
5P]BX@3>0K;4-]ee3+B(L(Q9+NB<gI@X3Z#Z4gcKPfg8X)L4/I^W[C.#N<3>8gX<
dcV#K[6J623C+Z8([RB,^=?]C5OB.Y=38<5de\<L^)e)bIR9I2\QCR3<,<bF(@0B
I,O]C=f5\Z8g\6^UD?SA1dCcNZX=eJbL>3[Vf-6TA3R0M]:5C5L<PF-UYC,/&DRV
7[f1JTM^G7)e\NY,1&CU5aA2JN<Sb4_T]\,/QQRP^+M^:D+a.G@->WQ?<LU6KT@d
G@?NMfV^efJPYBPfAX(AAa15b<=FCRd<;&)==f1^(#fgQ0E\<X7A9>U.:+P#?\Y.
+55[YF(JE,a7MYH3Pf>]XI^d[?EPILcX3C#C,S8UMVWSE5.GNVJ4SM4B1B2\=@ZN
P?._0?23:MZQNEePXd?>CeTF,82Ib(G[eGgVE9Ze8W12N1:&.M-)3UG?A8IZ^IeU
<6(#14P#::S,?VT;,LVdDHX0+;Ve67_<dNUR?I.>>@<)YG0A3BWHY970I50+62>&
Nc6>LC7H.X+UR3\EeUY0f.L9b\&7IEcfDc6/gPHDVHO3=eEK;cTG<@FbZ0DCAV^f
#:eZ09YaY76SI=+I42dJ-6c+<F_>/;_QU95\TXMXE.ZB_40;cT&G-_;1<97cc4eY
I2><@AG1MTRZc0J6_XF(-\WXd8&]c,@EfZa0],<OeAUAKUK[aAb3KfGLcZ.).W<<
>14cNS;6QX].CRY-B47\0HVc_;_D1D6@PU/=/4/T3B[:g20<6EE8Pa;9O6R1-8Jc
0RfD[[T^8@IWZFOC;_EXTLBGJ<LW,=C:D<b[GB;8a#LBaLUSF#^&IXAa2f_NV:/^
@:]S_f]Y=-3Q.I3KWE5[Pb4CVR[GPb_HT;3\9P6ZEHeEQ8W&cfg&2H<Y4CAYeYG]
3a\R_MPI0F]5<7a?4E^3,UCEdO4S>B1c+,GRSMX)H34?g.:B2/K8VSe51GF+N?92
JRSd;(a(A>@(J/<D7U&;LBE4<f<2ESZ-I.<VUV:ZPcP_Gg/4>U#bTFUVg/b+#7Z/
aA0f-^/X#HY)b<L@6BOJKB^?^EDBJ9]4\.ga3/_UKeJSBgeg)WSbfd3-0Ig^9S0M
.XM5O),XF(:/^HND1GH/U&\V)P8#X^Y;dWYU]Z-HHNS7g7L754CPH^P0X+f:f5DL
INS)[T?U>FVV95OaR>dgD5-:NcCeCPQ>K1<C]<bR=7UL3YZ/f,BTY_>[4C1ROTP1
f4+N/(J3e8/G<<8CT6Wg/&DP/C<?L4d.@N&DIUN1SH?0?Ngc.J6GeA/LD)fU)H(Z
E\dNOYAS1&Z\YgYAV3M0A-dX-;]ZAV>g,JRcGfc]P@^FF>fY;bI7N\X&,dF1?7E/
?8JTaUOe/(\XMPO_DL(b0U[/YFVT^]HV??CN1;X8/1b;CDM1.M&M,C/eGgMa]PCS
UC_a[:9X,7:JIBA1)1D&NV\9ZD2S99TP.QgP\g;E^E_P,[6V^548K1Sd?93^@+7E
a_bHHF-B[4ZS,AM?a1]K@M-8SAT#U5F?O27?D(Q^ACGSW:+5GK+)F7\POJ?;.#]U
@(#JAA^V0b)9280&&G_;PBHe@c.U6.^Rg7];.>IRF&76DJ(HgH,53&C64V2YH<Y(
E7VJf7g=0?U7#?f)1BR@MM5>6JVT.caM_UA.342O<bfC^6Jd=)68T^Ue7>Ya^b26
cG.JB6I=JTE&U5(=)38X8<0Z-Da76J;=J56)Za@4<>g9)>?FL2C4SbT+(^DHVLc8
Od##_Y=SdRW-?e>&IA^J[WK-KK&2S&^WGR1N/7I<>4VOS[a+d>I8EYbE)&U:Q8XY
XgN:gKZB.S/6B<3=M:)5=GQQ3MVW6MgLc6W)\4BFDa;:KRM+OP>_E34Q1&_,)b#f
dJUA?JD_7..M1/5=FPJ5LD@b7bIH5]Y,](RE0+5O\b782gO9?G-C,af0]VD5HE[N
C^N--NE#C+J^]W67(#3CE:)XWE:2(B5<=J,9\Sf\;KTNacAOeQDf4C@KX3dX(VBN
K/+QW#0_TdTCHCWNQ>,MVBbNZKA:Z2+Q2#gB11Y8-R326/c)_S>D?TX)-#If;e(P
&cB\2<VMDUH-D.DXeY>WKHF=OU1SW<JfLNG@F=N[A(TG/g3ECTK.:D9c1B9AAg(C
L+(0>)G@,4JKBg]8#:RYg?ZXW(&B[d?I.JE;I[NaHZb?+T1e?W/>@614C;I3(K:U
L405J[=XaVT>1P=+I:=BSBPDW&\a?MEIWXV?EFX-TaKX@#>BGPe8#O4c@f?^4&0:
L.>ERDJVKZN3/cQ.?YaSa1?eb17]c#fH@LBaF.ED&+Y:5U6?_9^#?NB&(TLd<bW0
41bN)#f])5d=>-3[F#)/YT<c/[6KRIa6AO,TIa=..SE-SUADH8Y]ON(@@eV66YR\
-9Y1W5M1#VVN+XY6(5;/H)B=,5ee;8DaeaY7LM:T+7;(D:83+aYQc5HC_@Ec]4/L
^\&5\-?QU8H8<>Jc/bOGKR?<CGA9#]4;=UR(F./D86\e9U7<U)C^E-CR&/<[+cRU
]V4)8eK0=1,dEBaW+3]MGI-g<?U-5g1R0<F;g[RIFdcL@-6WB[-25,MUV/_\>-NI
02T7[9?:ZeF2<Vb1X^PJ,9F5@<81L9bL,JE@>H.0Wd[#PD?KMT8Afc,@3^:YO8E4
SVf&dKaJSU<bOMRBZ4Of57<;27MZ<_;)^Ea1UA[U3BFM93[bQ^K8-#bgaKA&R27:
4bZOK&\HU)bMe#7fO8aTYe/8DJ-_BcYf+^g/^&,DF.aLJHYf(V+)Be;1NYSETX[4
L)S>^E^LE?0g7UeM5Q_LfTRZ^9baN]&B.PeT16YgQf?fN)JH+L?I[UARY5=O<Wc>
DXb^:JS[NQ(?I65YC4)N0[L)T35ENLg+O(_/Bg4d^6(#:+F84^6MZ^(LXZH)DY\-
daFP=KM-:g\f^_G#8UQTf^Z>T8aQQVOZ/2RRWSH[M5ff).aA&2MIETM&]C_(.ec\
DdT^Q-IC6]+,H65&?ZLR:6YDZ\)N1Og^WeXHC73H;2G0Z#-eFE+S0/0bg(c5(/1U
F>b.+)-X3)2Y)TXNQd&cMJTbb3e2_P0X_+9VJ_@R:2GU]/(BD.bbFT0\/M[d;O[Z
),KJX\HKZ[dYYNTa23#<11+:HH(SKVeWK_)Cb)>N;FX1D?W:-?6:<&Q8,0>NV(AA
<JUKC?/D?aGS6T73QbKeVOQXMW9RIOCOMGP-b&Rf](ZYA&A^C.-2T25J996V:XK3
V6dTM6SVYgeB4)@)FC&d/0\RJQ2K,;/LbWG:GO&fbN\=+)b;?_U.4T_Q?N.)bQg9
T+U:QZJJ07^c=);IWQe\=J/I^_:H?[a3TM8b)cLY1+4=bA8e-8X7UBBgUFXLBZOD
0XG&S\X]HOB//(T.\AR7g416:4@OFG:#1g9:T1Rd=?66)Ec&1/6U]F,b/f@&&/JG
A_2WQNIEDPE:&T7dIe>&VH+^cO>LRZ6K,9eK+^+I66K2Oda5Re&7N(JBKQdLK<gS
PYWUF4bW(#GA@T[?3,D]4_d0T_O?D7>5O=8Q^XV[4eVH_He7?@F-:M.:3=@DC/AN
6AXFd]SaS+>8g9OB1>baLaJV^8O:fSSKb(+V=5gS^Q[A#4EGBK^0b]4fPF#Ye1^Q
N@V942,#3BPFOfgQ^9M9;Kg;OYVJ6#?BTRB(8eIY3.8=fNR5N1K.Z>)+3B7/ZV3G
TZ\C[_)__?>GO]@g#RD@K#dd>OAEHV7ID2,)Z#KfO_\gMX2#M)0A;I39F#)dBRf1
D8[3(T9HP^bcb+,HPKI-X)(0;)fT\=T+,J#XPPGdLQ#<9QHO].T=IH)Z#80#MUQ,
7=#B+7&NX2RA7:2Gc&1NPL68Q&7B<W]U+KXX5_GI9baOe8?,IR14I(?NZ39NP1]T
UIOR=_EVYH+(=eVbc#[4F<7Ia0:P\Eg.V#5<5P1]Y:EY)OYeO#,e3.^EH9+4D:];
BYH::I?-OUA>_\EE<\(YdOS+CI9(.0@;.K<J>_R;c_@^XN+G8Z5WW]2_#[ITfOXZ
.g^O=<G>Cf=7W\5_=X<<S7_X4T>5QT<:add(B:+1dR=48X-:EY)8IBAbBY@&Rc,)
CQ.cZD(B&g39G4^c&5\4XB]4#J;Igd4FHc-5b=3L(D3O>VXUN/A#-H]Y_WAgIA?G
Z)E^DA9=UC,)@?a10^VeOH+UfU.E<_bV4M;g]EWdM0OG(5^1XMcDGBKe8Bc156U]
bM.LdN3OZO(KBTaK9:6(d<GcSJLNe4@Y8S)K^S.cIY&8dcG>F[8G.SR,)a\cReE3
ALA4:U@EdH_^@b4YB50&4+D9T=1ZVUR]3eE0@@(6N&A0aH2R^H-=a::/[[?E[T\7
ZD(Ogd_gML.=&E)7]>Q4?f/O:IO?.]d#:bM8gS3^G7M&@[3D<2R@B\ee;BDAR1LV
&=L-+IfE=PK2B?RDgYFXB99>LG.N8J3:1OZVQGaPLF/4Z##g[(NaE73N3B-aPZKS
AM7bR,WZ]Wa.W>@53JR45C\VQ?5KB2D]EdbQ&;SW(\,(1JNU4I<=U[1,7T#CW-g4
M5THY7>eO8K(:R+Ne3_/(BC1Q6dTI3=O++bFSB2S0O=6FVR,3cZ\g64,-BGQ#88d
-Sd(^43&60_5HgM,db3.GN#?]6I>N\=]Mf;4(B.T]SaQ.T@]ZSFg^fA6PM<[1\Wa
ST\/4@50X+_A2-gV:\d(UH]<^.fRS9D:F_?A8WePXAHK.gLUE,1L;@I9)O9:cRV-
,U=5P/WMA6FTMfXWde)P:P0F><eP((FEA5[HfDcQ6N=FTY2#57[?]fBY1FTQ3DK>
JEE;;#g3CC,F.]95&QPF=/WB)[0AfeOeNXZ1HKMUC\QXaE=BI?W-7;4GX^KG56V&
/XB.YS(KCL.J]CDD#EN+II\+\DLEa-Z_:-JEW=c@bM2B&)M#G<-,WZ(\<g:cD9(&
&VG4B-;&/fUF^DG6ZT;,&([^4^L+,0+^0+cc42EX]ga9JA/=>Lb6[P#XMfLIJgXb
&<aga=O<+(S;5+d,[<G]d0,2&?]3+DaT@edNQXXOCWNJRMe28VO<S:S8M&d+U>H7
;B^SX+<2.V#_)74JT@Z33I_42XN:QLcbY>@bT]W=5;5@4_a\G_3ZHQ?WFc&T,D.5
^S2>3?6G&Q\Lag5.,dfS\SJfZ]3HMIfR^.3R^0eD&86H\I(AF_OLISXJ;3EU6,f_
36)cZJf6-[SC-(Lfec+LM].E5@8g/]G-HGO-T]-E;_4O)d=WT(e]9F5V<O:gV1#B
7a6L7g]P/Sc\G-B#NeLM<26-Z9-&#5>OHM?/G:FO@;R#>HT8.OMYgF(f-U4APU]E
W<66:FdE(TQ#5?g;RDN:\=V[JDQ[D.^Kdd=MO1-?eV^a.b(X@Y4>bf9T3Z3bL=[U
Na=E2A^QOVOa[g5;1>NBR(c:bG-NcQ]HL_e<d>R82TWWAOV204VVc_\M#HJ:>5.d
3,..[MZVOdV@]>5Q4F;A;16V@L_eM&78M>M@R.R<[1&:.&3>(V26eZF9D0HJ,6]I
JQ<Vd.e.;>GD5gMG=@JRT<EKFS-N,I4I:[B1PK[<UUP],Re^:<^I;+&OFIe5A38>
d/5V1bQPPPA.VU>f)^N62-#V1D<9I#/YURK7,[4Y);_dfZ3+BAa8Z?4KZfVHKJ)&
GZ;#/VX\?Y+;6]LTc#K3JLaNYaJ0^d20B?>]4BDB3M-7M-;a-bA3:dN7CP;8;A,1
+<<U+/LC=^9]Y&M41#A>+a^U>Gf[RW8-#2K.GT>8JI=bA#>>Y@;O^GfgN8&-:D/Z
48Y=CH._/BI7Qce?>)[GbIPg@]fbBd?TE2CSZ183LcM^OX>CT)7D+.==/K4YX#RG
X9GG&D<5cRDT>1&R?QFY,U0#1=&aIT\2(e;gMU;CX\;c0,+]F,e_FIc<S/@XI>Vf
KW\-S.0V5C#Se]7\N[Sg][3^6gdPf.GU2:(a&XEW9;4,0&Q\eFHPNW:;)\Y.6D^#
>f+a9ROb9cPYe(59)GR<\6OKP03CX\/##bCYAIKVTNG=PW2V?<]Yf37YcFJV0/_e
(LKfU-aG5e2YUDO/f)e^U/#Q3D+AN/H<-00]I0a,ONb017&2A3:O6VT3@>E>\4/F
&Q,[c,7U4ZN?H3)C+#GC5Kbc:@fI6W5@EMQ2?D21/(LZe646L5bGO>NM?E@bI:O@
A.WaE=aZcF/QLJB]a8=@,7-XZ\O:2RA94DDX7>)=<&X#0#-b57UgJUTMO@8LF+e-
[D_Sg<5+LE@-GLdNOeH;A<Bg2D\.FD4RXfdb.P-?ZD3.JBO@CfX2IcJNR4&1C,A/
c+\a\Nd(A>B+g(UT/D]#(_@XS.;]BQ2V67Wfd/.RB2[,JgY&9aT(+fg;dTR;MYF]
cW4c9bKg+a<Pa:##4>c3DSUOR5dV2-8dF@EE1A\T6?_DR^F&2,XG;;A?4:KF(9-g
d2M6YQJ??.IeZ@131.E#:(:eGEDY/?UE4Vf#5Q2@>TW;BeK2R?.VIE,,2TXNKQ=@
QB.XAT=CU(A>eS5#;_g-9QY[R=6+;GG?-N9?6,A?#V/P1Y\/B&<X?KD//2_2cg=&
Ld#-K&)YQEJ>>[W(:K;f[dFV+BM(^MK8DXc,BcG&00?>Q-^3c,CG(.7U(MCH?UJJ
N)PV8#B5-\Q>VF7<Y&?+\L/;M<&fT1=(D)c1\XQE)GOR4UD#Ea@]&]YVUQ=Wd/8H
UEJZM1=d628(]E4ZQA(&>Q]F=WAKRLUF9T(06WFKcDLMLG)&C9B,C,e[R?Y-ZIg5
]#c=f/LAEaOTa&5]PKaM#I5O^OU&@#HY@4+,QB+85QWM,K7+A(RZ;Tf2G6OS>)P>
?6Z5UP,9+?d&8M17Gg3X(T(AK\@;c\P1b&P#Ka8BQ(g?a3@ND&3d[Q=6,WOXMRSJ
@0G7[P7d+KQ#\D],;:AR#F>8f65A2FPd\>PKJ<N:,,OJ9gCPC)5>b4_7AJ9Wfg)#
ST8HeJ:MLeeK>1YcF6J(TFC14fL5DOd5#@=]-NN-I7^6e2[6NaHET1bIZK;Cf9)?
4?\PDS8[9g702LB8QPcBRfFXI:UDIF,V[/&cO97._Y7PKE\J./&1;#a>0>F]:dc/
NC<Z_+0:;0Ef>]4I:T+JDTda5<;5B1BU;FIFbfSU;5@N_6;eUEf<8CRJTU=XNFVV
Ud,<S4NV#9J#-1f<I2-W:,a4X7&?eM23@+Rf)Q?E^H;K2.EEOLbYN5))Y?I1fccS
+C4&<XWM4;AQV7g^b[JK^3>U/_7:H:W4H[+T;d]=Q_-GT>N&b@1DBR-Td53KbXHJ
;FE#]0_egK&(6PMGPJ2LI7DdC_-K6_aQN(C)f&YY+[W??&9;+9]GK=P1[Id.RD1T
d5@J>TG.#P96R3OE2P@@0UX+19g2BZ1Q93/54.(?R&IEdF1L;4515G1.SH(-7#<#
E]PAZF-N4T&SH6-A)R?_KOff[WXD/D26N7K=bJQ/b/dH2>2A&)3D#f>4_Z6Q.;Kg
6G6W&8V_EXgg,.c\GIXMV/I:8QTN69.O/-3_OAMMg0Md&JYHcEe.^CODMcCQX.O,
dB=VO2T;2Q1AgNYDY[#/5-=HT3.?E[&5SS3\[8_@Cda#YRZQ#1&0DG\L5Aeb[W?Z
ITZQgT44eO;J;)T>,7WG3AVJ8V.^V(A;9V^gO/7?((9Sg=B@g/PgZ];7<DBHgU./
>dc#e+0U;N+L\Ed3>]>4GY;)X&@1EZ\#P-FYUM8:cNTIf?2^/#-g715X44TW=@+:
@BH)Wca)U61F:b_K)a8,_Y6g_W1/EFQD<.-#_/._A@0&,^4GMgQ>UHg>VA:0&DB5
NZ5I=KG[\0.6EMD/M^J3WI[bbJEUaOZ+;W\4C2?Q1=2Y_MKHF/8KJ1RJH4]\[MZb
5dL(aERXQG;\^77eYAbR1T_IS8+]_Y1GL[If)UB:G,_N_S61[,\G[IZZU>BU.0[;
N^.F4I1db>aP>OFW<L[[fTP#;.AE=+]8]c0]S197[a3Ja&?M+^+.):;cBO(;T16E
PMfHeL.N[.+R/9>I>/g-+[?.-G=R;IdX;KF2PD]ZPQ3@XA)((fEP#54PO;V.R@U+
R9T.LgSR;d>cS_gRd=NMDM<8&::GQXU<T6?4[TA[)+VHNM&N>3S=-be:X>=c?bdg
UPSS/+4(4A28/T8^CSg^Z.&.RP;8F4#8bdI0<Ufa\/HZ5T41G\.>+#.N+IMPA#CN
&UcXYI276?Z[UI\c4@UX(BH5I9)8<I+f=JZ_8eG3K<a-^(#R@/S1R]_G[S4APF:d
YU-G7cc4DUV,8K2@&<6[UMK8[T7>L+UMS[8S0F+1A/3g7)5]>P#ga6f:0d38F@DU
?]Zg>W#,D@4&\F^DN3Q&ZM9b39VS:@B7O:^9##d,CX/M]9EA9[V()2^+\>^Z<_/+
/TU@f_>>-2e:G>;2L.LE63&fFF-,fI@EB:)X7E_P@5;fDKLU2?AFHa37U;4#GDL<
KS@gBTPCM^8??e,+A0Y3IEQNT\-cC-,d[@DWV<P;[LbWabS82CJLFMJJJT5aXgZb
ES,=_HN4W;-:WJ@aTMS0/S_R@?b5]OZVI+_+DHaF\_2&6eQ4)S8YLN^:P:+/GHdL
K],TC[&A44BbUQX9&\DW#.>\PaJD0c7I>af7JMPNQ2P,Mce:g7)g_=6e:T0\GS9O
(TF<dCcbGWSda-<cFETQG/MU0T-bFYaX=YVRVFZQ\e@-:-&WE+N.]fd.LA\(].\B
2^A0c8-8D+0&?IgY+C/M/Je:K&:[^G_EAK70dCL315Y6Q1.3A_/XR)_MRJ9RP4Xf
H=c.8T]Me.H?2,cA02\PT1N,R7FT1>LWFZ_?_Ud&+YY.\VB+aEfT0g2K=Ob(D_)O
U=68gO<_F1@L><,-1>YKA,T-gDBE2LMK48fP1?<3J&VaDY:3,5R]1)-Jg_ULGeWB
C0WA0d?]J\&9Z&aNdVc#NQZ#B&aBR6?_?-2@S;\I^b]LO,b6.197\0.BcgI5RIUP
b>DMN<#W>W-S#;0N?GH)9S4?OIU&Zb7/KcOMOC89IYb/#]-NN,,U8NP&cB+07/H(
@P@W&EP7FAa1G[Vf5d&.&+][KP\83_7I\8c3LU;6TC=WW648:USA0>F#^]05@2MI
1,TWE7H;,b12Y/(99-G.T#8SdL[+POZ&cM46LW(L6;O&I<5K7?0M_::E8.<#:Yg:
]EUJ[D&&=<Z)XDIB]eJWV1^<CC\J-T]Z.9Ud,NTI_G9@KfF3X5WLS=>X[_gD2?-B
F(TQ<Wce,ZW;J_Oc+Z&-fL)ACD1\M0Z3-L3NI,,P[6eUM+G=Z)LMgY@C2/\I-Yg\
)#+8)D>KMB23:E6f,d_JO]PCgD2EN-ABYB6c@TO_X;RH<ZPHHdfIJ2e7O#.]V@D-
FE1J+9&)eWR30)IPFLB8=Mg<f\HU8d?/\]6-d\5UgQW29<YFBY72KYEL<3CR_#_4
G=(0HeY[IJ885.<-Q:;K554G(71Se?3-ILQ6E-NYB8f]=CMHc4<PPUKW=O9g:8?A
DYEb1fD/Y?+MdN0cE@CMdKeM#<UE7_QHP6PLfE(0V22g1(82dd#;eYe(c-,d@F1F
d5F3fdF+]ZP;LJG1<?OX&.VFUYJZ\FNLFK88U2A735C2I&MXW3;>D5Dd,K_eM421
TQ]1<?W_S;2QDN;@VQ;K]>/NedAST\;VJ=,+&NO1e7U@F]TFSWI1RL8Rf+D4D&g3
?d)7;4-1/MXIC>CGOUL\/dFI572?LB[_@<A>^5EK^-;7XNPA(B[SC=b<Q..22<c_
F,:=@D-NN^G^.Cd:4@T2G/bUVYc0/TPX1Z]G<I=SG(dC&fWP>?:cP4dX,fKU];J;
f./fNeY/B.KS#ZJa-@62B^-1W(0A.&)J3YZ;cVQ/7>Q;cS5XT=SA9bR<Y,2L1_K?
44-5\V7UHA2dF2=dW?>+R5XSIM+WK\a?K,W:Z/475d5Z,/2.K-7.H6#/YLNW/3F>
V38CeBQCg6^STR>WJZ69/,^?_Yc.P>_NcSL4>N&b1^Ka)IPfFaCQ7/7NO./<e>;B
@1W^BMdDGG]c_(LcY9>IL-+^Y)PQ)^.@1W-\[9AX;;g>XHRJB:e66D-Q]Sf5ME@+
3Z2DFY+V=8^VM,COGLa[>V1YA?\M0c-AH.-D.&dG?9Yb06T806d8(@>f=M4J:+(e
&FW):Fd=c,N^2EeJ/;GM7E<0>:CVb0f/-5-EH.c=0/P-M=Z_8cAQF7^#DIZ.(,&Y
,@=Nb(bQXA^,M;LY3BX]GNT.Hf<(F(f,,6\7+6/UQV:@+M8H8906ZJP3+6UXa\9V
7R=+<TCS98)2?9e1P\LO.X<)CH3V,cd@CHW;P./aMHcc]]6<I,A.O2>a9-EZWG+H
HG9YADdD<,?)Q0dGTA_NaN]T:YSY::L_TWR&HUgE+:CH^17C;GSe_&TdP6B9aM\6
aYU&Z8,:c>K1eUM17U=<.T/.NW1+1^@Z]G9g&<VPOH-,I<6VeGR]^G_@25/UBMQ>
++LP5NKdV5SBST3dL8]Yb^L&L-c01TY5HAZ_AL(RMSeMa;^E=TLQbT(f&0KX+&dc
+c68.]I(4I=UGceX/1>O=NaJ.CXc>1aXJ@@A++@K4WUS-ZQ2V5[1J3:FRaOaK)_N
J6e]^4&2#U31H#4VUcV-/JE8bSK6OO&ID9]:V<;c^Ic?09T?OL@=U^b,9)VS+RT5
eBH..<)[ON<EXUXEc)&.M((0e2/dZZZ-Z@Q5WNH+IR[:XbS2fD,_eSN2XI_;RPdH
C\IVJV(VDb>9b<fU3f?O8,aeKJ:9#X8P45b(X<32ZQS+>4S-fRZBU\/ZCENMUPRF
Wd.0eH8I#KAHRZZcgGT51gM16LeD;;2G3IY<VT]9YM.J.R8WR(MdH:VW=:D&SXd^
=fLTeN+5cS8TfYBa&WCW;\#Z+gF7f?KN9[&TFe)QbX(+MYeY/)63EbaYRdE=#:8E
)><EA^B9S+7^(8cVFdY&A,;:E0C>O0#;-J=RNVV=SP+VdVCF69WTFOX>b:=RfG@c
=;A\O)gWfe6)KT8=bfJWDV+/.)>4>_L)+A1L67Ia@VTXTgB(X\J]3bQX8d)8d2+g
^&_<73JFOc)S;F-L?Z8N(0UZ/I]A-K4BeZVA/bY2E&]&dAMg?4cUY2)aLCK19P@;
)8\X[LE:,84d1?<R3S_63FW1LQR+91\+S<b2+0ANW21AM@-dJ5-.8067EGHW;+75
FWFUIPdVU9+Z0J1#bP6/TPN,2=3:Z3EL6L77C\A:=b<?T6@IHX_+E;JJbUTC#^4c
6\3[DCc,Kf0.V,bCWgNbW8;#VN(&f>Y)1IQ@:Z>J3O\<KKL+.K8YG4YY@YE/_-f9
EVgS-;7^L)O40RUSP1XcPYK(W3-bERg?Zc<ZHLTA.#Q/C_0WC041NH11L4X-W^UL
d>T3L^_?K_YI:H:06eR05dTBG\d:N/CdK.dROKJEG=g^9g.TA28BS(?QBJK2UQUb
/D-1OQPBS927&<IZHf<AZSF]baQ?#4LC\TaU.U<Ef.#-A(Tg:XZ&SC\Y[fKbU>\2
U-1C;<@b[XNLK_6gC4]:R8EK;3YUH2(WO19;I/P\ISZE-T(R(b=?2:fUSE8ASJ-(
7H-^L1,OD93aMXd9V1NT3W4:DF]64^)9U,TH=->OaOZ]Df>E+AVD#4UJWE>#<17a
ESb?.U0XX<09N3FMF&NFc&.]9ccg(])A7?-U<]3-ME&cB]+^acCgGK[W&]QCDKNW
Mg1JMHS1f@4T]OOMGM)#adUSUK=gA4UW8#//O@)?cfX6<^.cA>P3MdD-:ef#;ULe
<3F6W&SJ^aM<-P^HbC9]EVaQJH=#MQ9NC#&ZfMgVHg3]7LGK6G?c00,>&1_IbG8B
5;DEB@:[QA):SNI7AI945f>JUd/TW[F7^e;/.(+/&=UJARVace6YG>T#OXe;>T;C
UcP93VC5Z(ZJULJB2?E6[>gS.QRG?=]E^H\B(GRWe7)ELX\LAIYU1]MAg6b<Q\[@
#[3)GEETDS=4>T/6B[VKb>=Ze9fW.&He3bg\KP/Ha-U7ZSQS._FM#P:&Zg#ZUF-0
PAb[LS#g#7AfCU5P)RT[OUf,2bG>KXd-02T3NI7&H3QH:+G]8Xa>M+?/E6I+5;79
9W\aJ0f9MCE[eT)@@S;AU?5A,FSCVBZ@.#:;:SJ(SD+c_A1CQC[8TeRD:JU3P<50
RF0(_PTc1>.P(^Jc0LeP8MG8aW3QT,Q_PMSYeXCg#Vd9S1\2A1X6<-<)>.A^4ZVU
ZfQL5M/NCV?PW]<bN6gbSEUQQY2/ED^#b&ZPVe64AgV544L02#fQ^5f9LdI);2Q#
OX_g?^W&9.7()cT,CBJ,@[<[F_\M.>4<B\Gc-N[-YQE[IUCL0&.(EM3_7LD(HU-]
Z,3Cd]AM@5MM-K-,.1U5>;^eNgAd8ZfRP2B8&3H;NB/F7a>;e7a4@B;ESC8;:P4d
7@>4.YEP(d:.D6=?28RY4E>;IH_f0GT]4<_;/C7a_JG9,^6CY5;99bc9)-TYC/=6
YSg?JOW94VD,gUgca.2)f;QH984R<)9<<5LPQaQ>Oc4Yba3<][X7DBQO#^U#.Ifc
d>^eP^Q9<Qc8Md+2ZG5Se7_\.GcW5F:Rag119>#UXD2YPH.d.<0C1<,aaeYJTeA[
S#,?\gK-_A;\aN3EDC.6d;N<+MgGUK\7366<RYdHH168]4H-9B^L_=4d;eO]<;8f
S,ELCc(91CA;fOSY7\._\2[VACB[XZ,XBd3R1.OUL9c6Y<AD;DgT=L1L0;YZg-O\
27@R.H2J^G5\g)+JR(+J(9&ag^VEI@,6K[@_JaH9Nf<^2Y<95/_#=c;LW)3P]TAA
Y;Ce0UUK+O4]AfKJTaT;#>R4NK2/b<#TeIb<b2Q]EX,:KeS<>40\:3\4?KWTEd63
#P9;+[gD]H^#BE+.d.[(:XOB2)21\M(f[\Q.<1,>c?.\f,([ND6,2/?Z9bO1>(ec
KCBJ05R#J=X(B6fbGUR8I8,a&27;D/Z-_7fG>@f5I0Cd0>&cY6Xd.MaH5\E]O2G-
=,JO#^<CHBe_)<HT]X-PP^e2CAT]EHZ=;ZeG&/;c;f6-1-]F2G&<8aJBDbRbLfdB
5=Q&L]F9<DTMYAQB_)=U4[2+P-(TX5FT7-HVX<&9[X8>^^AK-U_>eH-(LJMKZ@P6
B^?OYK?,/78ZfKR<O8b0AVI-O;,X[KC>(D;FD.Gb>63J7FW;KMN;Z8d6@P^0afF#
E[>dXacP-[1I1;fAWQURK3Z(ce>]<8@G6^Z&DCA1\F)<MER@Q^FRY0.@;2Sf[Y0I
5YQJZP5QYTL@BNc80^e;YB(c^KMa+1WfG<>N(?0F,EOV^eM>DAV:;aQU9c)(#dLd
[B@=VQ+[<<+K[<5e^P&B=I<7.@P7XdYIJbMQC<X+d>RDfEQY_X6V[dTg5V]a&7@Y
)(:/N3YP7,H=1c?Pf]]0G7)PNC7<Bg9AF)eFX5/OdSKF-^4NJ\^,eA&S+N-B-K61
-34G@1<1,Y,N9HW1.37Pb.,fH.]\U1],.@B[?SHG3W40DL0d_(0K2c=W5[8Z\]DV
R406O&5NDeBD+#]JTQ@=[&MAJb6Q48Ig(L?WQYQ6T2beWO<85?bF+bAD-@=fCWQ/
\6Q9d.P0g\JNb1?VB)^]X=e70a=G=+bC5W5\.Z>1,W94.AY0/_>D55A62FSO+16)
AT\HD3_+Y2IJeSN5A\<X9d3A-g1;K/>FQZef:.,)]DcU26CX12MUV<=.K(C2O5K\
D5#[ZST/.(,fVg7F]b#29\Q4#5PTG\I-f(SP^Z62\bL#=bKZ<Ug7H-N0S5f,[#\7
XKb&;A583c>86A(:_3]6L-<2(N-[VD9#WcRUK]TOeXZ@.NOeFW0(dBDe2^,e8NaK
-3Q(@M.L^>YDMZ@ZS.Ngd2S;,4LRQ.VAO>]>5:MbP&LOW-;db.:L-U>OZ-bBH/@A
.Ne^IP23NfAR\LUU8X^]K,O_\\>9&;0AJB)+Q#;dFR=?[32\NQ^,YSG2K6(C6#5a
H_-RI9#>eL@eI+>/Y;OHWN[-+]gP\A0^\R@,>\dN)K>M8gC>TM\?Pg0=^Ua>Yb_b
LO>@O0G=]_J/Bd40efCd7YZHQ&<4&=R;2.ZNN_KOE>cM8e:DX-@LIA=98XR0VFM_
5^;14137#&J5egbU_Ad>USK^E&DNf:WJCZ&+,I/7DN10K)Fa+CH>/=N\SC+1,FI/
T<Y)^.FTZeY[&T9\>>X.(P&#BV4Z-;024(f5db<bNJ\B&+[L(R@<bD=(f11J_4gL
^=X[,9_^ZGK;J-eRL?/Z-&JZ;S9F^FWd>[:S18>FT8dEaZZ[[JX\T+BbQg6[Rb4X
@ggBIDS+AB7Vc^JRb?3?^B3D21GG1X5HKZGT&WT<AYOc-E1_GC^],,[5<=RWK=T;
eMIE5_gg-O8E=MJ?OETI[#.[>QD9]-?SfV5AK^c&e>P7J+I^41MJUVW&[=&PUS8d
PTaRfG-OK20Fc(Z\M/B9XfMdU5QXQ7W[&=Fb5G8b4T,dI-<d0g8JabG0bLb#/.I=
2]FbZ<MB-c=/7_NSUT_\@BUEUP/^a\bZHQ+JF-KRG+OZWOLe9ADB(+K()ZFS^._.
ECOf?Q^BBX&C@?e-A./Y(#)D\#AFX01a(6[^=4P-,;B_4/O+8)aK?LdE1g21(P23
ZKEZ)a1&.7,@;QXY7g4CV>a,a,@6>0.;MF;Nd@D6fg0>]CgRcd]75)>.N+I^THf?
Z]7S7+I<6]^]J=;FAWda;F#d;-):S?KA9NK-c)?;@^7-O,<1K]Z#;.bFZ<.,>X1N
[F8MeIUadECd6>d0>ZQe?2QWCL,:],IE;S]e:>/;@-a0a)eB))1[d[RJ08I=ACbF
I(-@H#NLH[QAd^IW-_?DC)[94d-^Z,OWe@+/A00ZJ?70+KR[^Qd5AD]FfEfXKU4]
dB+9NB)bTAVZR3J^6FA2[dQY4TX0FCFdG<TY,[#;C1D7c^F<>b.:KRJdL/<H+FLD
[<WKXL-?Se1.5S&Y[?/G1Q/.^PL@geB0Ie-F1R?JIf=W(4GSAXM<_Pde8KA&U\/.
<PPMKQgXgA:22aXg)-0S5H#-JV@Va(G/>eR?G824,92<L&De:D4>0L[WPWeX>T#:
7EBK<-V-/I](Q+:5^R20cc&@HbT>NZggRTbDd_aL+4X-8aB@62/NI1Z5&We6Q82P
TC>7(/OLK#F:_Y6G.Z1eCZdcE4A0Ga;L)QgTd@BC?<bCWOB-HKJY+\(Q6-:@HS4\
a#QR32c;;PY2N[L\Z^F2b6^;,39DfS[39++6cI6B_51UAHHL7P9]#]4U_]Oe]=/e
^g?1/#f<?A+U[>N9RG>^XW^/^.OgQ2M@?KgG28K334V0NTL@;JJXUgZG0)A#[?d/
d2Q9_<F\/EJa2^1/S?;Kb[:1:N6fF/=2EPbV]R)8CSgG<X[X3>QL_fGd@+-=0P?X
>70PP9,;.5]67^)-J[CUN>&49SVV_cf;B.d=UG2[/Ya-\\<?fW(6_&Q;3C0=1_5T
bQL3?]ZK\[H48b]J>#[1N7d&G\f05aec\@BV=6,A3EL^O<A&,a3+(4^M#<BX[JIG
,c;U)BL^^:?8DVF0=3,V>Q8)+gG]S/67R:8X#d;fgG;Q)BG+ED&bBe(4YcK8V-E&
.6&QOe66JK=+6P:I5_TCGUH3_@aOH68MP\<@.S8(L3Y.2IG0^_bD>g_-(72[fOcN
:R>>\eM>.4aC_-(Z9^BB.QP/5?X89^<_f05B/Xb42:G,)Vdg9-NUgYcL4>-XGHbc
&\LO2K5ZSJX_?[g@L(Z\(D/4?5G6IE,Z.-]:g83FFZK^V0-12)U4K#WO#VI<8CP-
a^/P8X46dAJ5&,G\G2BZD,=M7fS(_FYZM<Ea>b]U9E^91@SX;RFE6,6=Y>8e.AKQ
[2@V#4071QYO<,W/T<P#8A7Q7d134fXV4H5(:G:?Te;KJ]^GY?9gRaUWgQDP^b4<
G::F8N=<_BDO[TIJWc)NT_+HE@@fGTNe,N#dIF@SU/@R5gN^gKS[6cbKLWO8D@g=
))?)&49>Og[Tc@,M3/GT<6<_=8CA@HK4I&^AS?59X8g/dbbI;LIH(gF,V2]ME<1M
\(_A.D4=]8TKW;OX=&/H=e9c+CWS_SKU.88_B.66]C=aN41eG>@J=L?b+#5IE2GD
(+=Z(4YMf<WBXX:RJ04O@D1eVI8a];9/:TV_V84e[R;#+]>9/11UMP_)9EW5#@IM
BK4eM;Z5;^/6Qg<^ecT^e^AY8_\B>ZL]+].G:4/0ZcDeef+=TE.#([:bG)>#Y?MU
91T,D7KP5T<&_d2,CV#<eXNQ/^#O>JPTC^b3;+8I6-+f@<\J<T3abWBW,#[[7Q4]
WS+)-CO3V#XA\E)BSM7=L0c8?)WN_P37cK=@I:Y?]F42RK8<g/().d+A]J9\+STb
f&/0&^b2QL<&.;JN[U)RP.0\e5QZ4SK_6c_)Dfge/A\_aFEEP-1?BC39a/+M\dgF
eZQF<)GWTUQQ\UDG>I6MZ=W5)#=(+aAYY@FY)-ZN@gf)]192Y:/KE)ZYU_KTO+Y>
/],AWSG.AO/KE>bU^)#GSdfWBDL=PEIZDaXR^S3F3D,@B],DLJ(&,;4c@c+VE((9
BHGL+Sb\#8aN5B&R;9^ff7]6RJc;LV][;.P^:DN:c1Y?0QbO+FcEf;,W&<<M2)S>
Lc9UYWPZU/b:JBF<9FEHI;V>9SL,JJLC6PXY7Y#J5Q\V&6[FREe?aeD<-/MR+6/#
5HJ-_C[\fSNMHe8=9fIce#UC[AAYb;9e5Y@7,f+58Ue(;/&<G?F:5DMdccOH=.cC
AWR(OV_XD\P<A=O1F_1g?Q+),-HL:B4QIb6_d2,SXTR20>=ND#)c]_W)CDSDgeF]
T,,J:NJ0.PN0RfTd+a8f=A:gTcS7TaP&VZ:^(bfOASF=@3H;]AEf)WL-ZS(cPg?c
Q+Y0e_03#:R(XMD4HO^OSB5P98)+QHEYUEMfSUE]2f4A8bKMc:-3:Fa+?MU2_U\1
&-YUQ#JWGJGgRFI.L2gF]._MD<&(&RMe:(SK)E/D&GK^KR<P:7.7,[GALXM)6LIF
UTME[\REIEF5ET=[O6XO;]-NgVNIU8;?C3[-_[\T390.J8/T.72e9=W(^BWX;@C=
CB6-0U@PZ^D&.>7X78I^:(eF2:/J\bg1,?#a.+7OOWPQMJ]XaUc(6;#W4/bSXV.)
C^VI@9fbT>AHf7@0Q1ZRTP4&]P)7PefdZE19UM-2F@Acg7M_(H0YU#C_@VMIdDN_
Sc6gJcVK<[Q\DDbXG,\9>6e-9H;G=GL@&8Z\73#L/f>IHPOaEJ8R.U(CU,>PgCYc
A][\Z#U6aP,QM=S?3?>L#)3Yc:.<I_NG815CB^f&8DG3=bLP<1=#YGU0LRX/G];W
#D/7b+\15#aFgYg(2),,4NST(5M@<D6:<54FA5S-AIBcUL5GT=bK77=I_=,aQfG-
H8C1+OU=,;F1#+gU;TZ(8]DD@5OdRf&MSYBe_7@,dI>7Sgd@bLfGH6+..(RQ9-WN
Qg8U._&f(Ab92@J;gYO_TSGP@Sa/J?AV/8<TX<M?eC\7L5FVH&H&N)GR<D;0?9Lf
L060],Rdd6+9HP38XS26Bd#O=<eJMT<P&-V2R#BeK.+:PPRAV1B^Z(7Jaa/H[@K=
]2OE]_878-IS-K0A5?+7TgH024.P96G?0ZX/(8W9b8G?><Q.RT&G/IO,+&;-ZMYI
:I=+J@O?H82Q+b@A4.9I&/[GZ)N9DL-9LM83\0&50af>OI4)/JcFg\EY&PSf)Cd0
ESc2I.2STA.Be5_dS92E+ZKC(S-BbFb[6/2c]gW?]3;G[NR1f;)LOXYJ>+F;A,)#
Nb&\ZWGO_=E,JO;7ece^3CC7^Q?9/]D6<g@[#>@R1.c0LgZ,.?R=/\GM++G2W4b(
9Q:ZP=K^3B5;d-Q-6:XIVPMH0@f9SCE3=JQ0G.;-AOd&.L53/d2c/a569[^gU^M(
6_D74[134L@R4#/G>Ef67SU6fXVb)#bKcYbOa979+R#C3HFWL1,</^fP]V?P9;cZ
0SHMDb3);8,75\5C3CA96&BN+;C9;>gPde:-[E)<H([HZLJSB>(19<ead#HR5OT5
I,PU9)#&B-4NA.eUY,>;27DZQ^)(OTX5+Lb5V4WR5>Zg_eRI+affSF[]dSf0,J#=
#6g7f2:R3\8_GH&G[S/e7+-)S_?CK7.+gT4,E:)a^>N(f#MMARC]d863M7P;TF?6
U5f6c&^Jc?5>CS()&7JC3TcY;,;d0OG+9^VRRM<+9#bGR?Z5[NI,D^U;3&;e#^\6
SULV>2MfPF+LFg9a3V:PD)-77]@5@71EAX0=33S16\^X^,E_?I)T8\Y=>=b4X0+,
@Y>828;d4PNP,EdV4V6.YM.)8)J:>C\E[d-[C4B=R.3a:1&)N/=Y-CD]0:6a4OeX
e,FW@T@U^.5TSI;MYV+;06@B,KN4,@,+Fb2J&CJ/]A+Z;^@F7^.WRGRJVIX1HWL7
S_/,+9dTSWVa=2]2ALXcV;[_:3aLZa^.1eZ6X[49[1^)()+\YSVfQPLU&W^+D6(V
T.Xc6&g7)2)[L2gLJU&F55]c]N_JeSe]+P8G0AC01KW79SB\U^afJ4Z/55&#/&aS
DKOgX9.R;4+X9S1/_Y[8M/[[,=X.@M[SL9?>2GZI8SXXIA<Wg0(c.][fEge8cF+I
cEffDOOP,GdR\JL-aW\1<9RDLJ_g-5^-C+_0J,HL<4-FAcb<LO2I#dE,Cb3ID\YB
#BFb8M4ATH-:,f_J,1WNE83Of2Q3>F5WFE/<V/<[2\Bb>-,0XKWN,X@3PB:L\6[-
N.U651(;EUB+3<FR+4;d8SFOB2>G=_>,TA6N.16cWA#JO=F#)7UM/PD[E[VI[aJ?
8AKfdLFKQH(/5&<+6OY4:G=VF&R<\?^D07.d3NH:_H5:L5\ff6/5(&TGGSF81e>]
EPXNfGS5)\afO,NZIb?3#ce:L&#8c5F4@,F=bN79PS=/F.@c9[LFW<(>L&=<W^ZK
b(,>;Q8N?a1FIWW<^MCX>Ef1/KF[NUNd=:I?/(AD.BAP=4R)6>3/1JF:W8]Z9)RZ
WbZfb_7dT.WA/N80Ta^7WKP(ES5A(NIG,/VU72V2;PIGCEB/BWZH:_,VDB7S(P8A
+J7A._Q&JN-7([ZEY?LSTaE^UMb-O#JGCS]@L8?;cJ_:I9DQ2SMc#UX_gG4.,&O@
C_4bZDKW7.2(LVI5HS)b913OJbX12a2)S4=YW3&Z8[V)ZM@L:^cdga\[.@GX@^14
T1FD<[]II3Q-A??GJ3##cg_JZUQSQD/G]BLH[RD,b@Vf.DfMVUOYIC(D3X\WY63?
32Oe08eP\;<WTN5FPVDIe.]Y+3V=4f\:f+VBdQAgFC=OYZ5[.<#(4dOHE-dVM7VD
PW]+8)H[K/bM03)9K@2G)2T4GD6-/MCDN6F@;_GS,gLX9T+J:Ze?=V+0RFH19=6I
OQZTNbCG><a-e9JI@3fC7E5a_QN54MWND(C:#>5EO?gB\U38IAb;_HH6:+fT=cZM
:U4H;RWNM6#^4\A4L=U@()#ZXA:WaA7b)<P^D4d.Y+eP6e[>LE;E^P(SS>M2^^:6
1N^]V30;.O55R<3HE=YTMHZf<H])_=_[_ZB7A^-V0Hc])Z(,XA#Qc3Y,.?\0<4.D
EMgT&#ZVRTSE6d)<MWCD4DMG+8X1E@ec[TT2Yg9L>QAR/L5_<2<F?W;c[#K[D5_d
,+>UeK<87R-:)Q7#P#Y=IF[]aJUa[F^.g\>;_NQ3/CAV6;L^.e8EWX&Mf4+9?>FO
GQB:12Zbf9>F1/7AY1PQ,FHCXG)L:W[OfY82VX=CQWCAZ5P1\d<QM6HAQI,]]e)E
@T62-b-dZ\Fd/-;N4d?RX/DI[3)K9>Hd3e\^&NLcVR\:SX.4I[1]b-Rda>J)G#,5
8P81a/5c8A+B5We8DUYT(9FJWdVONO6/#-990g<bF7g>#,d.SO22+N4VC8M)Y3LH
,]26OW9K@E;:D^bgPWSN<dBXL\(8O5=L;P\gc8fVK@FVYPX11QNfGcJEJIF[eJZK
#I+DXI(-/;S1C-W.F:B1ZaW@a8,-+Mg_+6@Se\)..Y=ROE:g<[Y5XFX,KgP:<L)P
3Q+QBKa=daAQ3?,-UGI:B#;.HY_)3H6WK[)Oe0L+DMFTBZ9:T0B6:gJ^Y21>e,Ob
-0H<^Y)LM^J=:0X,Wf^eZ3^P6[X=WR_2F9V=LT\S,Hg+X?RCWc-\efNPWNQI&JOT
GB+QTUBBY53:H9I20GPe:UGP5TOZgNA?P<136)@RQM-P4O@+cDJGacUV/JJ1<4=\
H:]T^1CG=?PWLH@.,]CEcXAb;ICVe4^?SZ<3Ca1]->L[=QaZ,UgFc5bJ,B)3@X[]
?O6WKUZDe5)6@VW>4]+ZSV:I6Qc8T63f5?)]^0Mcd3>SP97B+C4UbI6_5F8IJ=Z2
/\#6aAS0ZOXIULUC+K9KcQ1_NVOc+)Z:VC&^a3KZ9_A0,-P0K,.EcKHPe_1a?AKM
g3Eg>C<bS-:V9<Z(^V6DFH5HeSb2LQ03IdVI;YJALJdNJF<KX>F]b8N+gRd,X7V^
K+.97+,e)d5TIc:LSNE_R#\WbYMDL<d.aMc(I3+LU8/VCEXg3RKYb=3fI1_&^#E)
,BW>E/<Sd#M?O^^-+::38U5)0bD4:+A_:GJ2S]NIM]6WSG+UGGN16]CRd9+@[P38
(.M#(_Q69g,c]/V.aU3M_#7?<,>(YEf07@^4V6KGR8Bca,?CR(GEO8RKEHgK5KG,
WBO+N>Rb.CdYNDQL\<,E#Ye#N)R[+FWfVDT,Id,L4Jacc?LNRAbeIdLP2WMb57W\
NSKXIFZ.[VL@;4C#CT3;fDR.=JDfND/b#^00H2,>:>AIMYGUKZD/cSYD\F/FRUE6
>CX[21&a<ae#Xe^LPLL2S^UO?QS,P:EISN3^U&]])::WYAfEPVSAJd)e15?7,DZR
O6)O]I7L4XdgU-HWa)-.NZ3A8-9GI3UPPJ4I?c(Hb[I6G.],5B9HS.XNY&FX/49E
?VAN&MC5dHP[](:CA5B?DLId(I>_/43E;=/D2)O]g:,KOMf8C;Te1dd(/^I)DgTQ
<DP_#Q)_bQFR+.@gf3g>WdB;\2OH7J<+<DT[BXDY6g=O2>[76[4[H3>;D&c7-TFK
0_/OO_)>&BbC-TN\3ccc=gD=O<Z+1Vc/MO?6&ca\(d_g;@N:AUcC(<cdE\aI0.]5
V_f6R(&Ya6IPaHC(JHC@08JLa;Z9Z^IZb(&#76(\5RUB3D8VMF<XMXIgVV4eDeA@
1_<,T)@DH0O5E7U;D19H-4<Hd1V#O4dJK;^3-@g&6d>Je?&.L9ZG.gROD>U6VFU:
LeW7;?CQe,\dAOcNZ_JZ0Ua7R+B,.G#ZNQY2?d]M3)=>\aZU/^?<7@^X8C7PeM2G
f19R/+?cf],FT?8.?K2J3,^Y2VRS3A;S:\B=))dN\)@e=@1bg0ZgGOCa+9N85J<2
&S27GB;K7F.&((G2:G5d=b&-;5UMUc9UA5P]4b8<6[#I-E.dd11&Hc&28XA34FEG
Tg>1A@11G8_/6OHTIOC.N#F.KM+S\47eDg:=#>&JHHLd].@U8EB../3^R_3_4:81
:#N^&a^((;SFAfW7S#>)MMIR&<=R[?-Vf^d2JcIFYX@/38)NOg-],^T?W_>g3c,P
VJJHaG1]3[cOZC1IKR6cNCQ5A\QLf\C^f(M>[VQ[():V/7GU5V#dVXP3,WDabJ]O
RNB8D6KU64?YSA:<FCCK.C;@5AV:/HMgb2B_XIHJe2G/e&6a)I]AYA;7LGVJQVDP
J3X?Le^W7g,X17,49=#<R?T?fQLAT8(b_YVcESY?+SMHI16IEITWW^aE_?EZX0cL
C7G_[Xb9@KNP8N6WQ].MYZO)^8B5]c&db+N:9IP(1DWM>W5fg4/);KLZ9+DJCKW]
7BJD,VF<@<f(;KUI.&8GZ#bC1d-.;PCWCK;^-TZ1e?BS0\[(Ac?S.C:gfM8W]1BZ
4I4C+X1J<K_.S<P+D1(_\<]DdZ0[L,F;YDCH&>b(+J52ZX=5\;S0FCL5;KE-#^JF
+#5O)K@.D,0gO(CaT6gRX6BRB/^3<49(MDA00R-ZLZd#WRI<&CF)A7S74Q7S&W5f
XE5C+X+#=OX^Y@_&]a,.QQ?YCX_+;PZ=I?>Y(:?P@5L\#ZE12G8YV>Y,=A=<g2>g
Zb_7P_>UUc.\I->1e9_TURf=aaRM&YNBW.,Eg@H[Q04SNWT4Z?Y>.,A,f#O<(4(W
2c]g3Y+I,S)3YGVC\)N+;@2<YfMf^JMNH++[U;+BBU-&VC1PHZ3?MX^X59fDL^XR
f58KA)V4gaLX>e6.Lb;9+7QOVfO>]C8N17[2OF0U)O1d4HDYJS/e^A=)&+@,5=[\
Y.)57<+D>b-(+^O@0A,VVO]),7a=A4PIGcA=E\=d=C^.3X@=+f91HUP)U&)Z_9#S
A1A@(8c9LU0GGOc8S<cG[+[Q?B6?SXgfY7X[==/1:c1J4Y4M,DAS#;&YYL>fSLNA
X2P)O>[d5GAFe1E=\>SS-ITdOdVZbR]4@+HX[DPX?<[L>a39I]M,1fVV>?_6dPX-
NT:dg_TH\,4C1ISQ),OC6&9+2RBA1+G@B2W3a+G4EAI:.L/FBI;J\F[TQ-.8gIWa
FZ?N[7PM2a<SKGLbU>8L57+)aACf3-egBZPIDF#,.#BGVTd>2=6ZREIU^Z\<bBN?
bE@XfUTd1YMJeeOIC9G0M<-@92@==UNMA62LO^7K]eg[7:,ffc0;GX45>;AUO1SB
M\CXG(4/0&K,bY\2dU=0eFBZBZa(@(>MCLa2_g#+6]/2GONbY.D<>#I_/4JP:7RO
#P\+c[MS-=ICRDIAD[NNH;8=CJKYMH/+7V\a8Ya>e#NN(DZ53W(VP49ED-bE035M
.C\;[(VI0]\>Kg=91Z74U=V7J^8&<\:D?0YXP+T[91gJOQ#CY2eFSg(M/VU/RU9e
1VC<-d_E(4HE-51(eL-eL)(0b;aOS+PYKcRCB@F4_)NVW5dH#NW3I7:Q[&W.1QWW
@^N4\>W2K@Nd4IV9AEde;H-#_DR_4Z#8Sae+;N-1R1Ng>Q76@VXg/AU@0P:J8;<c
YW3aO(CfX(?/XJZCgUP2Y?O9/^Jb)^)YE3[D-58W[DLgI8gLVG?TL/Z6?AAFN1CK
N+L.KFE<^(N+2N.5S;C)dUTG-KC9SFFWVX3W@9EV,/0./+8_<Q=(;CSa8)A83^;M
FE_aA\L9GLg9S0(5>SINVFP&IaQU-6<U8e._^dLaK4I/?VRKegg+1&P/O=B=>^,4
AgEGF;cH)7D:fa,gdLK(-:d[LTND?;/GU&c5D^NF4d;IEM=P?&dSb@<;Y)Tb62D0
YNZU<3LaR3J+^+Z:H).IdWW25KeS+)+dWf+\G1#OTO0N<P_/_V\28JaY/:G1cC1e
=X;QHE_K=SV:@ZO2WL>:(^GZJ27=dL5YM:eST)US/b-:X)N[E(Y7@X]3M8O06ZOX
C8KK8@Rb)e^=P51QBc937BEOcdUR;(MUVL\9JNd-)SeUWZed5R4U0a^:LcTfGHbL
YFff@P]++d#.M8cR</VAF74Y0.;U_BMS8F[-Fd^<ILER6;VB09gMQZWG^O+EWVcd
9^^(/P,-BD]75+\F_&J@;#@=Bb=631KB0F\&cQM6WUW1QYQ\dRK8bAFD/1Z.U#E[
NBY:L&YIH#Z2>f(Y^P;PWSUHR(g3&=\=U[ES6P:c#CH2TY)43?XYVDRO>0HIaMM=
X;<]9DdZ,3GcIQ)Nb#HA]GPKgIT<3#5^V0,QEBH0@TBe\,c4c@[W,_^?P.K3(6bW
ODNTJLAP(2d6/DZ0g.#+XEbPIaE+V-gK5La??43N>)_J5OLf>G#-JRS7a+\J.[JW
4#(8JDeNCa:6?FMK@B/D-C&F\K.O+,c>[<bZ8/^N:3Sb#8\NBffM,?8gaB3N2U@f
TXddDV@[0?3CS8_CG[[LFd88VEI=^]NH)b-gF+45?0-g:2_.@L62QR^H0eJe,P^C
.H58A5<WP5]G_CPgf5SIRF@+M]fW>FQ_&</dCI7&CCY8dU4DX4]cT5KK:98(T\A9
b-Zb8N)]4G#[P2/-Id=.OO0M4.^(B+[(WgMH(YR>NK>__-&0#X?f3g)-J/]:S+cD
X+(8(=5DM_W?09dF8B^ac?F>J>[6OePM\aC5)A-<a)62TKTcT(Gc_Yf6)VGRI1;O
=gG-NR45?6)=IC_8cCPc;BGBd9ad-Q?@+#OFHD8NbYe9g3(V#WBN17[ETH[C0&e:
W>RC(fL#gVcbRE47LK3YHg=#/NW:HG(#@K2=S>Y6+WUTN;YV7)L\_:2JP]J+[2/e
PPa_f,)cVZ65&L<g1F-+L6X7-\bd+gdPWYYH@d+2b/QV:8NEeFZ/Dg[SB1>H@aSH
:I,D1?[]NVE3[a6fIKL\f>9F:EJegK:PB8KASG2[>89Z=M;R.O6&(MW1Z3+ZA[Ae
:P+FL6?bLG.FG5&[TH:fcK_5>=B_5\,QXO#Z0V=,D[_54baFG6)?JI-?)Z?_D_B2
NI<f@[?fUaV:T,-Y__fNUY)8FV3#cU6PYEc(U31KUP?EF@R4VL][51>9YUJV\>&)
<a:3)U>?=a9T8+MBdFR]>DI;)AHMBE@T76^=Q@9_/\,Xa(5]8H(1E]N,K@[;E5K[
93aK/3F9A^J=+-)GbV_aHTKUNdgXUCF<U:/L+:1NWa)=@ID.J@__3EP[VY5(N]F>
1[/X3[V@74)#PEYAV[2(Yc&C3H9;Hb[.b^K[&f[0VZ8GDM\[=XHKOGccKDS:PSE7
Z)I0#CA0F/#1?46P&[[f8c.@.9H^T=D;e.LAXM4NQc&7K;<[b]<;Q2H-88];]72\
0;ULF1>P\QMY/HYb><\gZ)ZXKb4AB/OUeCUgC#eaM8C;,[gf1+J#(U7KN,&EGQ.>
6L=J,/N&62HMY)NfZdMP0U5CBRJ7<)M^(#L3cVN?OAQ9-7+6)d4J]EL6^-(2PFJG
F#_\gag>C)9HS3f#dZKDAT-[SbHE6)NdeOJSbYMdIeG)gP8U/McfNN)KgOT_aa]Z
;dNCL59GCM+TI8gB[Pff9d8?HTMS>B=[L1;H9/AE&//S>MTg_??KO)7W(Af:A@H,
V95dfFK3[d,VPJ7NC7L52)Pa@4M8JI0>bHR(JXGG1D1LCZ[=>bZd)@XI6@74Qf+A
NG-\Q:9#+L\<MAfA;.<B3N)C1X<W=,g8+T.U=H,4b13L/2#5]4M=ZW9.ESDReB-K
_CGO#6;2-AAQ2c:D6?RQdHH#GBW5L\535g6+HKJfMLC=Og;@.V3,C[MAeY/[IRd<
&2G&/K:XLYE<Z/-b5^N;40:c>g=HOPU9C25((WQD/G<J[V(XED)2;\4]TA.4fHXW
SPY@X]KZ8OXASQ-:BM7(DgSM);e(Q32&\]Vg[D\b-9Q_JY_:=+6gaeG6RTe9G2eT
FU;dMBe-V/0EO]+0aBH(XAeR[#c@]]QPS&\,B2[#\@+g#Pde/_KA7Kbe]BV#3d>0
H.DVI@R35;1M]<A+_Q:/J]<EE7/(@<f;a]V@@YXJf=U=[ebDdDO2c(<WO_8fL]Nc
HQT7I_I\W3<\+0QdS@1^Pf\;NPB-f.:JdKN(KJ3#5g103W5W;>H[@_4Z#I3CCZG\
\[-E0Z]aRHGH9?N947VY_TW?&^AC/6\T9a5RN\,_cb[,Cd(K6<8FH#+0#H+aG92g
M>aM#>J&E:+VK6P+,M&Med.]EU.]\T=8]^+0AWS]5OD07&S/@:b@@,UHZ^13@JbC
JDRV)g7;4X^17WFEHf,Eec+TH(#3<@Q@3Q\8\e#a\\32d&WI@@MZ(ZLI.e(+JIZK
c5A-f:2:9U/ALfZQEaI-8cISe2f^_-e1JEQ,;2HHJCZX[VQ#OaWD7CYCM,PH5&J:
BDCT.E/=a5,1^.4LZXf4YN5Ac(IQZR]6[KG;;Ld>c3^OSb<I>;+KYJX5757Y:ZJ9
AZXa]XDFNXW2QN&J+bOFd2c#DGdK&4BdJbLd500/RT3R_YO,W,E9_M4=JY9?40(A
:GI.9RH:G3c\>&JW/ODYI=FZ/_,gefRLNWNSL.(4[CL;dSH17cWb49g;f?K\WIYO
7G3=E01f/DWT<Q4>W#V4&-IW;Q_[1N;]D)F@RID>Y-CGY0+JW,A=F[627=+73Ze@
/YTX-DIbCe;g-1@_5Ic.UDETB4eTQ2+FVI1MZ(CE5G/^6I7Z,AQBRIB:IHYdPG6(
V:2W/TP/+S=X#+F[/<BYCME3Y2W_.\9,b#>_SM@&NZ2XQ.Ld+@Q+b<&(,^bKWPGC
e]74Z0dR-LVF^Q8=FeB=&9IPMgE+9([fQYeDRI,?[gS@V_.G6(_HJDOY7&^BVXc6
?43YDS;,U8^>gPT\08WdS88Z#+]6^SFX,[4T4RLKZcbK4=-,cE>2CU>(EJd6b]V_
W\Ee/5X8J#Vb5D/+3^&DLPD[>9a,=)GB<ZbY+-@gd:Y[6VE[AYU1]cd0M8[c@K>D
1.)?.bSNL&F-T7;?VbIdYLfGNQG6L9O-g3P1N\+6NPU:e;NV+]L:8EM?4PENTbL&
b7Qg^g](=0Qf2a(EJ1-BT2F>aG&A+=Q-d:7Y7eK&E=MeY=ZJSX)]-,ca&ZaQ4=??
&\a9RGV=5JXS0>Q,ZA8C,M0[\D>J>;5EYB82QW+6cFC1b]=.HX9#Pfa05Vae/7O_
8A):(&8\(C,)6X[:BcJbg9)bS_MeY#OG.)CTUg<d&>9WJM10H_.?HdP(=Q+U_QBU
<CX14OY-UV-&?6Z1]A1ZgH9S-?>P=>?S4;aS5f-JRJL]K8&aU:6I&,5<P2>&X,^S
\LQ)ZHR9HY9TTW4,Tee_3_f&;Q-^/dXc<d,CcPQT5B.M>&I.O,K9eS&0eV=R)V8G
><bc+[S<e7L@B,7+RZP-efKRT)<Edg\Z<>]6T(MR2@0TZ;+OU&bW[_S2GaX=I(XR
89[UZeLD^KdcKQHO>#D;9)WHYD&-FLBDb&G9EP,X+UOXBMe2)[<(4fT+Ub3?[,;=
K8bHWa,]b_ROKX#0cC/aJZ\J9dWd5_K346X/;]eN4agI7BYFL[Q:U(:,\+X3WZQX
DBX^HX]4_A;-,\JeN8Fd-;<A7-Vd>2(.;&J=/5^^DEd[Q/=cR.bY#RBfMW.7W&M4
-0f/[Jc<48&?REYSKGQY6GCf12O9\O;P&>LYPV,R5-a][6BH::2J=H2SU5XPKf;N
RPPFcT;?T[);WOcQT>F,=&GeB0Ee8H7?NM;LCNES:R1U/65ZUWf9#0,78;R<75^.
D82E91:.-03eVff]W8M=T)TUIK#&^#GRVHXEZ9]SCR^O8C(LP?gec3\M2)_d521b
GY.8ZgJbLaQT+>7GZC9[&g@f(OBR1N\Nb^,]=^O0F<06<UD;>LVY2aH-fLH@8K--
(Y.R;P/-W+T8W@dA7F6fS0@,eI4O\77C4L21U?1/fR+gbf+#DFS>A(]O/fZ.>X?_
M7gb+[)DdXXI\/OIe@ZTGB@\_8c\6V^a1SE]OdU2c-[(&f>/-A_I6K0:D1.0IeJH
QFgZ2]4B+;(,CSI/;F@Ja@dF<EZ1]RGH(.RTXDeSZN3&Mc78U[/]+Fg+JUT1@RZI
_[TNeDL2g:SC#;MKAW(_+5^ba+(;786RJ3d5OObP^^9/fHfG5/SLYRN5H>7&7e&e
OJdIeK2F:_dd]??\GceJa4dSD)54/UY>LKbY6f1@VJR1/S.1?R]E]73?BCE-CK@f
fQ&2YXP7H3=#V8f^.Eg<66N1;R-.QBU-4IT-@[;4/AgS0,=-?H4Q&a#RA@PSN^:F
;;M)Y\UD9-R^&JSQ_)=_RC8O3?L2;5?<3K.gCFQXDa>96/^/:;:0F.G)C[RAOK\N
9\U0W5f=@40DH680]#Vg\_:WHc0SHDO#4.^PZ<\PQ->[MA);E?XMZFD;f&EReELb
T],FIREZRBK(EJa^3^:P?.<<N-WC=BV[3U&.)7E-\\.cdT-DGfE\E:[Z;3/,ABdd
dg1c^YS/=b[)=B\&GHFHBMXU39a0)JIRS4@LQ]YH.b&)gRgJT=8.,9@c^@6\;g&9
<GSO3;dG>F&&;S\H=7F>Fd^??1KR[KJc?S.NLSINS[d8L?1f+A_/d2N(.A2LC1]]
86b)NeGegb&C)g=><W=MFKQ/:gUM<>D-1e9&QZSR15=DIB;cQ2JSUDP>^O69OI[Q
A0Db^A1-OLAcY><(4Y8fG6;5f&C4<]9F?T9.UQ<FcAeCa6WbEC,/[>-B/,[L_W(2
:SCD\(/,FJI=>:Y_/WbO6\SOL;:bWd4a2YP8?87+U=ZH<F]7/RALf;cIC_<14bS/
E9(5Uefab4cF.URG6^D8BM&<SN8Nb\;DIR,QRR9@1_2L0?FOFBCPS.Y3(&<^LH/G
G?0LZ5H8GD8HZ.;ZA5;4+(,>)JXZ_)+5BAc1<S-N\&EA,eH421\(If@E^I[+d^V]
M-B&9M:+\VK4_AQ[-MO[WPfY7Qec(dLg27SNL_4N6GZaUX-G7=+LS42,#_^dMP5f
BD-RH][^b:+eAg4IZH?[VCON>Od6?5e[6S;;\:8g&ID5+<WM)JgNFcE9g>(>4,W;
I5>3OYD:@+=\0RRJQ:Qc=7=cJ;>gV\MYO)HN7<#<^80E;B,NbCR7W0(&VCE]9P>Z
V533cNMP;\_=5,#gHc6W^(63ZD]@,L5JCQM(N9=J/#C\6H=4D;c]X1(@)63NAf7&
]d/P6,(GI\b^\0SaO?4.]4;L14YB7O6?Ce?RX5#G7W]Y,3L08L;@g]Ze0a)Z)?5(
B-@S:]C]fBA/]P=N3/Q@CUS[g_5JI,G^:V,3II/@8V5)UQ(5=ES+VSFT]WBHM9SA
/^b,ZAO):W/S8_6DGVUS;#O=>@T\1_=1I^1dPJQYL@Da@#P[^)ULY#cf</=-,X/&
CKGQ5K.EKcMZJSVNT]b.0WLXJ12.eR:PF<(K&&H4HKe7<IT6L>ZK/ML@4@),&bEV
-_X>]W),/:S2<.9SgJSS78Y-eTQ_1]KdM<K6;A2_GWdb^W\Q[S6XTQdVZHI(BMWZ
G36]\D[GGB<MNbPD(8HIJ2YI).g38>g,eC&](Z^A1,\GNLMWO[TR3PDRI;+;9e4>
9McM8P4SgA[XO,#K.S#KA+)G@QI-,@G?<gZaV#R7caSEX=NQ:ICHFQdSG8UF+FUN
6##WNO]YQeT3N^N)C4WR/e&C].4PM>WCQ(dQ#(&O0R8<70Ic_2VUOTaaK@K8MUcV
\EbX,W2G2bHC<.WSS/7#A)0B_Q2O-,(aF/P&#XF45b:B?f?DPTRDEa8KEQ)H-Q=S
E-]X6I<QA=9?a=M(;6^fJ8dWWAOUJE?DRCVVNFFIY<3BN.A^BG161?\>&D&#=5&0
#HXM1E-;)WgReVLR_ee<2]2NM]0GINeEc8Z/a831d(b5S(PgfC&RLM02GP<.dIdQ
J-DZAdBNF>VSP\?Fe_Dea1\P,@Rd),e2LQ-Q#L\4_Bg_2e_8BS(6Z2(.SOYgM\Le
P?VZbb[MVXZ.)1c1;\9JB,QM>55D]1PaZZUQ064UCG&g-[Kc0)#]_4a1?+/4gM\V
G&C19[([GR&,a>#\8^,MO8^<U7_U2cZ[#5a289ISIP9]e9BQK#f#T^g0+3cc)\O:
G1K&-6e(cP4.LT+Ab/A_M)FE58X>Of3B<ML\O(K1#-X6?&IMV4<&Z5@:>E^04O\_
PJX_@1(Y0H-G(1E>eBVOJ<11>7H>1cCN3c=\,PYX;VI5CM#.3UT@MR8>)g1RaG7\
I9B4(M[)=6>JO77bMa3@b;D5PRW-E53U)dSe/&)[T=R:>?eOUNC7g,<>&5HK:&@(
)XD=65TW[IUE[b_\),H?8)8d\(Og/RK?.fW_M4_9YaN>A<[[^a8cJ)aA)b/P?5+@
J.F+B<;-0D=(RLE?KQG,4&8P@P_I3e7];Ab),WG>EX<IK\XFfE6R?3,[K;]5[:C6
UCaDG?gOLY6C)HMB?V<bK1/FW_6EN_0@=eEC2R7ZLUDR8=Ib2XV(eJBF0YZ1ASb9
3E\GcFX6ME,gQ3]?e\8=[<UMQ?g<AKY(#6Sb6Tc[Lb^-]])&6eRF.X+dH=\T5SS5
?-g:<YN>cS9/\TJedT[J2@)@]b?@_09(8d40+XA>OO:<X8<8;Q-J<H,JC&,I10(6
c@X8&=H0W4dPHR#_E67U[2Ed(RIEZ008+ba,?X_NS=^Z\9YSG18CS>3bgeC4DB>Q
XF\O@c8C77)S8/S5g((c&I3CcIZP]K,8>@>S8e@5_UP3:8ba0Bg[V:XJ(8B]G-eU
_Eb?H5HZAZS(f6>@I;_Af0[D+\f)Xf/+VM#7?\B;agJET8/;+Bd)#bUf(IVMb7bL
^bXC<eVb0W<GS2;C01;I4&/(I0P5CgGD,B;B=<9/><JPOWd=>,[IV4R98AWeZ9J(
,CHO:-A4W[IE]-V0Pc\_8W4dPC:0c39VgYCL(b+&1=G7AD4CcV\5=L;MMKa0]H\d
]#DOK49M:ZOX>APN0FQACIb40FdH6(fB1b>8:9aN3U?UALAWF0:@aC+:L&Q,ETUT
TV:>)/W#7E2VAZYG,8dI5BOX(FVN9?,AQ[#f=>gA\1^_.2:0),2\[f>H+[ZCFUH@
>4WT=Q=fUTJJO4b8IZ>bL]Od#K)ENf,],38H5<b0Y6#51>]3T(4NDM^PaL=F_g]d
&A)&ZLJ(F]\J8Y>[=4M)#(Y-5(HC6[9P_HM/1feXK27[>f/I\UG)Q#5Kb#V^0]\&
E9IA.a,a?A19GSR\S(SP1CGIA#^)NR+8?RS4[D&X8ad3X/M#29g,0YgGc#T^RW/:
Qg/b15ZI,CZRB&VW592D;U>E)d#@/+:GO=g3&50W@50f[MNcX_V_TKS0H0O?BLVQ
1ON^Y)R&b5/RV1/869/.66/fVb<UQCBe]0:.VRQ))38RaY-H<K/FM.1OBOCQNIPV
V]IXX>f84<J&WU+)Kb7T_^PM&>?++\DPUAMS7ed=3YbBd0eJ<\VTUMGC4ac9O-SB
V1).\O=]=_g[XE0bHPWFSX#dQ[Cg#?bO;GI9Sc8M\(/BOcOZ-f_:O;DKDR@GVRgX
J8M/P=HC;53WTZ</#:UL_-g<J9+Z]-#7D_6O-HZ4_KRLPEB4DZGI<,BYWGY-<WdZ
SXT#Yd/8CW8H@?Jc0P]a/B>>(NH3OOLV8YM<<R[a?O]RZ]5FENO0E>@;+?6;c#WV
3@C?VHPK57Z)MI65B1a,])YZZA)EE6=5U_B#3Bg.7aG,XPN&;CO/Ag6#3(gSL3Rf
3?XQ9cb&UKO/G&Hb-_.T?3.2-Y_g:JLR6BV,1X6ea<+HN-bX7]]2U?@#?8+=JZcH
K=7+O::&K<QX<;YgIdPC;0@P2-IT/EW-JBX2bR=?RV_g81JP)LMQ-=OFfJHe_aQ@
((7B4^WSAR.PK/N&@R).,7cULUGg[SJWDUg2U\WF.cbH7?Y2<^aU6;7Hc:;1&e<X
R;WUWI/d_I<b=>+HWffSAM7T.A_.,H3R?71:](15If6XKb24:IHB&]FK;]efNG>+
ORTbb4)#(O;6=?RTZA;>W57Y+[=NJY4DZ48X3\g:?7CeT>[ObO,b-0[VO+7&^3@D
fNBU0T.XA5D0fHR3[dZ;KaW[?Y9]ND<V+,1)X_F:BedCY]<V0Z=^QA0)X)<5ZL+G
/\3L;dIC3<>#2A7H9DS6F9cK_S]OGHVK<@?\&]S=8F>HO&OH?Mb@B_3dfA;8F7Zf
2XW9>/2#K:\H4N/Y^;\I\=S0c&F[J-?,_H;Y#bD7>Nc-3B?5]G12^0]Xe\EWB>9<
DSUWAX)Zc5(V6Jd\9-A\K:ZBY9EZB2-VP.DSK;&0;@-BMS?A>,Y(Be5XGEOQbB\C
_6<R);&BA[&9O=PVK96,H@H>4Wa?(8M-0G10Eg)NNI&W(C,@18JW0O6L5g-J]_KY
_O?<H3d]27ebJ>5F&VgAPV,^4e42\G6_KUe4?)bYWM.T+J2=eW09UJ2A(P5C=0;F
;\SSGO[K1C181ebW[P#TDC\?TPC_E7S>>C]N=_(BM&_H33gQ;]X,T3QdEU+.[ERL
@(&Z/efcc&=#7@#_T#TH,>c(6M_R2MFae8A<_YB/;McLZ#XMM++M#RGdcbd[AF=W
fB3^FJ9Y5.c&Q29[c]GJ]=6/0:_>@Mb..T>GTD;QYCB(:/KGJETNJ]U@T7BI^7M,
,1f8V0CV2RE];_)0>Z_DB3LQ(S#\EU)]>,5J6WL:=fS0MO<1R)1Nfa-S]2JP,FC]
;f0S:/M>4^OIQ(FJ5R,H^;C\V\^+/>H\Z9<9@FWA7eP0,aea-I<>GdK,1+-V,P8]
>@TJXS-d;ae7M3+(TTFPKa44S=7\:LGC^,PGK9RP94EW11>GRSc<f?6-.IWEM9:J
SOSC&T\?D&.64AUVWCPP1aaO#0N6c=>Q1G>CKJcXW=)8f&f\?:M.7ZT.50J1f?^T
&gE7Q5(F+X2B?XQ312,67D-bgV3?AY1WJ6B0[RYaA_HD]>3;a5&^]Q-d>UR[]-\;
=87)b(AG3Hg70a9/e0g/4L&<a3<>@Ecd4?OZ^^RR1f?VIF])++DR74b4=dMCYcV,
9ffT.cI3=e.K/NG71?^>;^>#;E\<fJ6(TRV@:U7IZRCXFGHRQ0\:Z[c#^K/4/bG4
7=IU0BMa(7#NCg23/UG6e<5N&M43dE6;()Y45Ef?9&M,N&5Zc#;MP1fgX));D&L.
NCDC4_BXZCAfV1g>YPd8M[+NOHLUI(<cZ1SL7:1W,@ZU(9I^Y+FRT/@1dcOfb/@>
Z?8?T4Q88E29J>QfAQ+PCag5b/6HeFQ/#OH5II@GfKb4+JQ2;D9\5L63W?[HdKSe
-FOH?=Y<4Mga^L1I?/J1E+)VcXbV8cKZd;0B[A^]f2-?TH_@0/>&LG;#7f82bT1e
@F=cB<be=##T#3BOE&;Z/FM+[@AR+RHF]_^4MUc_8O,PN,3W0F5Z?Q0Z=WV/?=ea
MD/L&2Scgd&B^Zf?SJM.A<7eX06TeOg:_NQQO)/J@PW;O&(IY.1U9b(:56b.K7<b
CHdH];S_CQAIg=bJU/UTF5[-KbX2K\X8?=QA@.[Af1C3]f7e90Ea0VGDXfQSK0:g
\e^@?)OQb_ZC=3Q06SOY\80CBbZg?[12RP@fB-&?BWX[[_Y(^EJJBdR3C.40YY@Y
TCS@:BK@K2&Y0S(K4>G]A0#S+-=D5d+,8MWJf/3E//-6[XCK,,QMZ6P^GK+/K:#B
GC4Ue=bL;ULV^B_=6A([fSS456TYA5VND78FRT9USR?6KBcI&?C>2Qg2QE3=>&RZ
V#a]S6Hc2V2cTbf]^IHIefEXg[KBG))]a&0\EVRZD:V0bCZA>F@3?PD]R-@2.1dE
U07?4(;F2a)QQa/7B.U;.W,Z2(P_DNXX.)K4\7>E<KJbd0A^VB#=3e<LU\(,4E0<
QcV+9V2Ca/R=.B62cI<)MecZ_PN72B6-W[9IRc=,ZY]BJ5I&@7c=BbKca9K5VX-]
U<RIFd<e+&\=0XX<BUISb93:&1[SIVBM,I#.C7&LZZ(@/N#0,cY)O:+;WJ>Y.P1.
aA,[C79?7HG&C//B8>AZ,V>3a,TD[0fcEFBA/\8:Kg)R]U_E80M6:Y54O0#SCSN8
&>?EJJdbXK5-D^G8/=L@c6^cdCYK7c.OQ.;/Y=ZH28PGI=ESfQGR;IIG&<a79.E_
XC#_75M/7#F?Qb#PfKJeVJO_<+M0=dYM)+a8YMSDg\:K@&AVZ.AX9Idc>37g(@Y/
CBJB\3C:=W/:8O4^4<\VWS>F8E_fEBYAfNK[NX[N_bE[?V<6YXLYc6&A)ZObNc7T
3I^5dZ?ULT+([.+(D#/]H3RBJ:ZIARa9#C3gX>V_fWEDg-K^(T+H=1fY4OPR/]D_
\g0WJXgQ.Q:_TEZW>Y>X+:(?G[RaW==]\b>KM=cP@#Y;D3\\>30PR&aL)ZA(5;N0
7O4IBRVI2RVATDM0cF:?2FDUH(4,R_TG,<MXfWV_ML2d)+(c&WGPS;)LK-F9T542
,UN,O0^=?5T+#\[AY2Z?+SFG#XA/R]E0\RON\93[)=&WL+J4]D_(U<1[2_ddSbfQ
,1#1N0_bUBC4//N.2fJ(6TGgb]3e_K?,W_^YYJC3.6Q]]W&Ad=R@TC(IdcG1OcRJ
6Lb+8]Yf6aa6f0X&(^BR2]e3+g:Yb@GZKO[CE-&]T9(;I97#_B(^J]#V@]DTL@Ua
8OZEfS-?H)KH3b.XF^TIaDI:2O>77;dI^Y-^CVA-#-2D5)VVL3Vf?bD9TU.N?M00
441G4GW>6F[Q^5[Oa(3SG#4@>/]\VgU;c^KfX7ROB)[635GQW)+\cc0\bG81Q782
]C<C(4b-2>)YTGHM[K;g<8\3DIdS5K#OL_dCV+EfD4?#OB\9c\>\aNPS2O@22)eA
Yg,=N^E/(G@6D^PfT.aX]S>H40dA@0TY;;:THD.;N,FUa7&>&gb;NT,909:ee3G:
X?W3K(5)--cB\TT_)7/BD)].6eELYO4P+Z;81)VfR</2FH@G+^T,fH3SXJ-_&H&[
La8?^5V_9g0XYDK4ZN-TNR,>a+/\FC8_>3Ga\&O)5D+#9R(VR0N]HSG84PM5U+bd
0H]-?SF45>97PZJ0g3VR^b^H>5P\=-I4:eS8La;+E=@,cX)+[J05:F(ZSac:>QaQ
ARA/6<5bD7W@;<&dM0fS;,><,0JQVMbOP/JZcRbI[N3_9e7N52L)NU)3);+1)TZg
6d_K4)/G52?M@eedB3b73OKRedBL5HWe[a]U[JWL=1T5TCD[OQY9J:/,Y\;X<F-g
TMeb(eA\@V,URBZNOdJ0\9__[A<DA)bUa?)3,A99B=JK2+A?_N0<XTKd]YVX,I9S
c\fQ].JK^faZJ5#Vd9SG_@K;S84[H5;)eRb=PESabYB45LBBYT#Ud<QXadOJf,4<
2gd0/@KS<dVFc]^E\5CgWadFeM5NIb,EJBeBJ4b6Z8CDLP4e5[M(7;af:>U/DIZ(
N;,_^8fI3.XS8FY6:gUAMR5N-F[b[RLF)e2=Y_ITQPL88;fD94^Y.=JP9N=]-&bP
e)BC\>T75E_/WGaVMZOJRI/MZ-EgP(-#;CRLROK83I>>3ZQP?M.SZ=_E#ZT0;DN.
Z-H,eXQQR46X464XXL8eN0?@,4F5W:b08EF[>,LJgCCJZdd;Q4J)9LU>Z8CD:.CV
=e@_Z>gK:JI:^caE1I0_G<EcIf0<Y5=7e(^H)Pd-5=25413C,/ZdO60ZKO3f1ALJ
<?TFa@-<fc3Y/ORNcW30)-_R4>4TPP15CTQJg08+RS:^I/@H#&,8e0IBWLfFK5L<
8cb/C1##;VVS@/14gZIP9+J<<A(;=]\NFEVdNLW\b2@R?2-e5A.-7Q7BD(cDe[R<
U@bOKY[f4MWQKW(,E&8])P/;?@;ZA?NNG=.QRYR?/ZJegad\B@)X,c5f0>7;PTT7
ZV5RZe/:Y+&X/LAJAX=K)X6Z[^BECBec6E3@KQ]LK<f&<+H@?2I3L(@M8#Z?9VK9
0#8W9RPJPY+CN)5GSCB;CEfC,Jb,FfFFQIW?L9T9HSIeeI::Z#217;Bg97VGD?_M
Vg@OK;GC25&SS?,8M_9I2(^=2X/Z6XZG8M+fLS.#:L#P_<fCE59a/7NC((XEXL1]
.8E:BR9e);32PHfG_cX03CS7?d8WQ1,fZ.NV_7T1:A,?X5&e3D7XB@,dF)N7U0O<
d1/gcEST]O@81PV&C(+M9FA<aT,(14YZ@bH.\E3b+@BU>MV3:LK9]+_MP[B2M;WE
5GH&XJ&c[b0[S<=90H2Q>Q5_)^^>E&#>D5FgWPYHQ]7SKB+3+g8\fURA4HQKIc)2
bT510F(F7P06RaQ_([P:aFFJBCCDQW0?59OR[gGG-7(TC-VIG5,AU@^.EQY:Je;7
2COdK[F=3A_T+1QL<T,Y)_Y)/IH/N,B2CZdVI[3ZE+O:V/.N9=2a/XTX#g<Yg<#T
RDNK\0[,B-8Cag24gDF]c]750aL8HDY7L+0V,?)>;N_Q&X1>N>,[HC2S?H@>UaaN
TRYH7Y6MI#>HZ56=U9-=X.\3\6.:.J:\g:F@5PN++WJ1JfSac)\+G.@,1PGOUFSH
X&bE.5YaJ5=[-^/40^.b-Z+\K_06WXL,&NKYg.:4&Y<<NLe:?IaZ,L7EHX(3B+&;
LJFP1R_Q_;Q8QP&3DH9S-fG7PS+a-TP-C,=gCA3/ecZCG[dbdLW&b50P>.L/RTR1
7[DBAHA8\@_D<MKSCg.bY=JCMBOdY<C-?6fGKJH3(,FLV(M]@cM_HK+ScV68I]K)
F2,D]I,VO\BXb,bXQ7eQ.J3D-;GK5SE]=D:58(02AN+X(J.f8SXd#K,ZSGgaX@V&
8OM5Z0&\c0L9RH#U[f@Yg&O;YPGKVN<?b^]fQ1I;#>FCF2g>IRc&XSgM=JSJ:Z1U
B53G-^Qc3?H/=:.@?6D^E)fb4NN?-KcL\OBUDI^_2^;DcWa#]<Ugee\Ig&)c9<0.
7C=WDF4C53a^H+f^CC>UgSK4W,83<=d&M=KFYTRa_I&egV]U_17=02UL\G2PSGJ<
GO^6AeX-;PCF8(,E=H@]+3,]G:\Ne(,@@L_QKf9T1R7A[(+f347f5X:>M;^4Ya_K
RdJU,Kb)BAPaV=6;12IJ0WgIg2Z?>F9S.Z?VCJA]V]^PK&#d=@c1]9\@;gF7VfQR
\8f?]]U@G9/]2>C;g,,4Jd@^^W@X[WF_.S)gUSb8CT.bR38-e4Q[2(0L]1@K6428
^ENI0-?/Y^D2=F..R5/EMXQN-c8#SI>V1WdMYJSP7NJ4\Y;-KJcF8489+d,JSP-Q
@XQfRGDO8E:5R;/K_6Q8KI.7ed(0OFX=9X_<@L;9Oa0OC+-0d-a83+&TOV1P&J71
CL49Y?aL=_Vf2E+64cPRccaa#GF@;T8U.T0b;LdUeP?H1cc<O18QC-[RXT/IY5QY
@,F.RXW:C:T_E#1X/X]g5H\8JM=[([@CR=a)fGXX>X:(3R:K\XPY8B#[VE=c\2NW
gDO^ZML17F<7#R(TX(883L7BKVCLe;HUT^KNQf3E+ZCR_T5H\KL(VTfN1=W3MUgg
-dgd-K8XZ88f:e7cES2.5C_a(NN-L6Lac-D0G4&HDJJPfcKE79bg,.#cR60PT2S@
9BD>&gB220-U;T&;7>XE7M@Y33;e4If\\#0BHdc:c)29J32,H-+8[W26,WUdL;)@
#52@GfA0T,\d05NB<AJ,W[:a48K@gUI0=R0A[8Aaf?(4MWSV0CF9^Wb)3FcHN]M/
O,dDT^3fE,4+FPVaIBacG;DSVCO1FWDFB&4PR5IP1]@AFT9CabJ>QP74);>?^F(J
ZGeX:TI@#2=eK?EXW8XJ<M>BL]I0_.5a:_Z8gZAV[)\E.GSgG?S)Q<);?0TQGB1.
5E;WBE3O=U=OfH_3.[SaU6<bLVaW0XGYc=+Eg9-3<<;.-bRG1UVbR9PN?J^^>H1.
E_0.^c<RP#-R/[Z\UM91=A7W1=S]e0cW_#B/UYg4/D7R>68(L7)R^1V.>-GZDEdN
e,-RfX(3QY-2XZ><6(AcgW9<gP+JT,>37C)+G_[SM8YJP4;[W\8>Y19MU3_Z^0SF
Q.?0&9XM-JU]?N:,&SRS]OGE>Y)?P^3a4D\8T(7B>880PF9HZS2+<e/GF,NPG]6Y
T=JO9#?)2_0Fg<TWK9&,M?P@dg4g_4g_=L<:Y@d3Q9gQ22U@gKF\]GT?4WIg<H5M
B=SfMD:0<=-);N+BTSH:-32+W:^4,8Be8?g1\E]0J.fMC-VBJ5<J.&b#E-f6]f@J
<),-<6,MD,?M_SI-Dce)<TJagE_SJa-FY9Rb6BWM.()JD23RI8Y-/[9UR,Z\32WS
S8+X>GDRePH0ge=MA\&2&US]Nf,IN;7O>[^&9\8]CPWFC@9YZgHGJ]d8HF0@-D6C
+BeK4P6N#4/3;8\QY-ARFMN44.Q1.,I7fc2Mc2a[]KWb+]/92N1ZA:cF9bN].AX?
>OAI99EV+0L<aB7#;1G<22DS77g_Z;>)8F0[]XeE:;S,\1F:cP:T\TE5#E=UL/=W
GR0G/A=_HU(@)dBI8<[(=,HYMIR35Pg+ZaV/(_;#N:JVAK\H=P5<;P_&;,4,B?QC
e?X:0>O&[+3f6O6V,Mf,_6f<2eB7K)dAYVN&JM7W;;c8?fFD=N6XY&GX=d9,Cg=H
^@W7ga4XAMZ55]QGMc-#dbf4ROc)97Z=Paf;g\@<Eb-]N3#UP,&.gfU>,K(G\Da5
ANX0H8HB@4@^.FB2b:160EeAM&0^A6=VW^\A/R84A4#7Fa)N#/,^9;Z,[1E0MBM1
Q,#(#@4NDdG].eBF7RH[:c+^MfU<5J+[CM^=LR>E+9J9DP26eC+J#Y#<-./-,fKZ
UTS=:5;V2_<0BO+_76P+XZR@,VO;VK)[Ygdd^Cf,PE5O\b\LDQ2eZ74/N1@beI9S
BFfK@<H0;B.AY1.2:-YRPNA8,+<9K25G1ZB0R2eDZGeSB)c-^UEZ_-OY)_(7NgB[
P4^\16<>4EEcM#::[_O\K(?E6EWR>KT)-J:bH,C7d>E;H53I=LU&I(^H#eCca5eC
L2)OM;7F(KS;(7&gP-HbeR4,LW<f/66dBV31c4>:KM:8S&]C)8fe(=Y]XDU&O9,8
/Dd&FXO18IRQ=98fJ#.cF)NW9OK@J=_,76Fca14)?;UTQERL]8,5@Y;GX4Z@BQRE
][aEAX(<S)RZ<&KGSHZHX:[JaEWTR;@3O2LZN<>NMXR=9\DO.cZ_d4eTKERd@aJa
,Mc:,WcS(_>\.0,SAKd9IT]\)PdMLZAR)d+&C^(F]7U?]eA3NO-MN](FXZ>gW,e4
N_DPPGGJa>2f/_&E)-C4[Ve8C?_6V9UOVf?RMA^#O;DD=D61I78cG]TC&ER3>SO>
;[b2efBTR1#50?N=1(.R@FSC<9fcX/4eEe=Uc4M[faSf.,LKWZD<c>bZ2W7,7-J\
32aO1Ve2AN&=]:PWZeK[7[D#J@7b#)F5VB2T7<P13ddS/0@0Z69g<I7c-<-2QIXF
29\#:OAEgb5XWA/V:bR<B)_,18.PRbbJNHCYY&5-GIG\+.dO\R>\V1:[1AFd:.AO
HfdZ/)[e??^?MH[6:74NJ0/;/J23T(XfJ]<AK6f\[;[C5b;>KPbFdf;RZWXJ2^+c
XCG?>?D9(B2]bbF?)EA]J2@6F,WPU;gY\Q/N82J_4^MQ]bY;8.B.E.[f]V;A>2IJ
SC78&D^X07LL]CdKR/VT?C,\1CG5&#4./6EWZ9]1\^g2F7.N)+[OQ#NbRd2P+RFN
P(#84dT<>HHe>dG8_@>WgGASVQUT:R#V[@]^&L-&P:N+0P]-A.GP4K^TSN]@/,0,
Q,Yf?>GbZ&f+c8;A=#1(MN/Y.\TTNM.agS3#L95?]/.].MUW18A2gBR+;]NKL(5G
JT\J9dK-JD?\SZ=OR0]O>CFUA43LN?[<0OM2P]WG==2We-(M2.)/YXNZ92SMI(Ge
+K(-e#.\J;>T#S92?3)>S0_::RJEOIeCLdPV/_fXd[++C0D:5E(bCYNCI[7N/0Z6
PA9dU[c[\+;]RZf#9B^9]6ef1PI(WZ8;.@-\9?R86&dOf#>#-]+-<cP+E/K1)=?0
(b5<KM@0F8.CVAW)GAY2?d,1_^/e_]9AdIeE^UH[Hf)V8IGN^@9gceecHT\DB0Kg
1I/MFEL=@8>X^&aE1-B?LC[)@3(8\1c8<W6[e=A6^B^KIVdTW^CCUa2)A1bIJ<PZ
/LM-&)14[U&\H8DQ.EZY53;>R7[deY)T://f@JAB\8KVe4])EGY+4-GFY#dV;O,K
ML8@GP;S_]e3#IK0e_C#@:4g8:cVVKff>(7J9699Y3B<_391Jf[@PeKCc;7I<>dP
Z5VRPSD&:#(+d+fWcHJ7)T9GYB3#CZWT34,,ZD_RcY;gS]RSI;)N6O/gT/LLR4X[
KG_N@2LQ(Q>7+Y6HA05B+D6UacMQ6O3d6BY;Z+_8(6U6.bJX[4O_\C8\2_d,:N7X
dX;K<RQ8QX;X4C[)G4(Z280U,;WKI\\d13R6&RZE<3#H2SDCEW,C;,:dNfP_J[,2
2921(X>5CZ_SUTS99-1L7f(6f+9Kf5g2-6J1UAg&U8C-2G2@^Ib\g5._S+bP9KZ+
#G>e_(4cY??K7,[ebe7#E\S0)Y>e5P<U\^P.7Ke:c;NIeB]M2B4@dMFb38^[BO;=
;-cAX;5Vc>1WL7L>@#P<.OD8bJA+R;)IJ3c7f.eK@+HNB&:Q(^f:J@:b&M<775&&
-1Y<#[(fYEVU]2D-bgCUSe,a6#YQPS-V&M&gB_;+MeKLO9/7CT@2QV+??HQ:]8[\
5NAOe]2aCfXLacJe,=KBf_4+S2?ge:)P<e?YCHG92c<)G#AQK,>[;AABfO2E_b)V
40)@4f\>GZ01-fZ-P33QUO-8[,^2f&;;3F<#33Xa_3BW2eE:Of]^eV^^F1J&ggT4
2Y>M=ERW+[7Y4;FM6S[ZF#1-G0#AGOXdLYdaMF\SKND>=)cJbF^Q>Y/T)U^+XSLJ
[CF:4(<D[+2[?(&be@G?T>VeYgSJ)IeH\K]HIcQ-:;_Ac0aT.#5EEI]Gb=+8X.74
&[7F?d>J:@&;1dL6Vc:?__Id=37=8_;??S#83\?WE/_6TgGCZ835,FG-<I]:JDF@
60^4=IKf&7:ZGVTM@U&g8cQH/=gGQ?:_C6IQZ1BSI#;(2d[]B;IK/VD06OJ+[N<6
1#E@QAZ4:]fM<:/9dF+QKgd/>P#MFJ<EI\Df<.QOIZH?\T6@GLE74UUCaJ&+V4\X
]5^7,6.D^C<0b.e)M8cdWDC\3.IWEMU_>TW\2?]e..L^3ZL[7MHG4IW,&Q_aH4)>
]QH/R19_3H,<>:</7PI.CPA3-,LR9P/)/dSNId<3dE/MA^4g9<I]#L++(R>7d>UL
f9JY#&3H)dT^BSSJ^7ZR>8::ZEB_9J5da.1)PT:_=ZI1V7d86TARJD:M)@fM3g31
JS>\(]F#JFL4;::>5NT5H\RB1XAge,Q\.N-Qb1D6>^Q?78Hc8F8TZ4:MN$
`endprotected
endmodule