//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2024 Fall
//   Lab05 Exercise		: Template Matching with Image Processing
//   Author     		: Bang-Yuan Xiao (xuan95732@gmail.com)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.v
//   Module Name : PATTERN
//   Release version : V1.0 (Release Date: 2024-08)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`ifdef RTL
    `define CYCLE_TIME 20.0
`endif
`ifdef GATE
    `define CYCLE_TIME 20.0
`endif
`ifdef POST
    `define CYCLE_TIME 20.0
`endif

`define PATNUM      100
`define SETNUM      8
`define SEED        86
`define VALUE_LIMIT 256

module PATTERN
`protected
YU;NHM)&Md^U:?g:U<@&gX,CN(IQcMS>VKA35K?L)08^)fOT56P;))TBHQgZ;RW^
)+4)[=Q-3GE9)[IEPATcE#N((,dXW;4A=_Z3N584,0;Z>AZ=VUY[g>#?9e<99H?L
Td3VB9A]/B@RA/,&A<&HOX[I;4T\d._BQ[V:dX;@=Z)c5c[.1:;^4e7Pc,6U;;f-
2gZIebZea,YH-4Rd/IO0b5bc,-9d583;#>E,HROY&:67<3H\,:/HPYBK@9@<63+-
/?T;RJ9TLES6([YbBES^1>5HUJ^1/.27F7-U\&K.aZgR6fZ&3VIS)^SAa1C>bXY+
)cUPX@9-9Dg88XZEXKYY/<N)11I;.19+W]-@c-)eS<GDK5\A3P(?Z,JF.(\)5W3B
,4V@C(AO),B(c/HGQ\GE:5.[U0@:@Ob56ZTW_A_O_[9VgDB>)E?;;<83@JM-1K\3
=fQ2M#]>O<E)DbPaB_KNZVcCFc8<F7K7eE3BJ]AW>DOD7IT>LbMXe^07VUAZ2ZdX
XJ>47g?1SVMY[1CV.O:\F7,KN7,OQ5I=S&2F7A_>\]&WGFPPJBAQ634GR17I4-KA
H=d;HbTDD7M6X[EL<a#]ITK1d=;<W2S.8BA]SI&^GZ.,[L:[AD9Y@\T?+[@:3KF>
@GQc5NWEE_fdQ[aL/G5MY^CFF(Z]XS=/XCE@X\:Z(?LfKL.9&Z3WL)]ZUS@bD9?Q
-@;^.g=S#NPP4UM^RLQZ<T>CQO:,0MT=86W2-PJ<a&X)Ga.@&DCW8((0Ua;:cTCD
TRR0D^LMEH0@_&PFRTY,W]D/):;CdU<3J<c,\7/H5E5K63(;YEDJGL6[KHX:1R6e
>9I3K)NX+3cC0/L?C/dZ@M.U3ZZYT49gIUW@L,@-=+<H(b.3P(0,-RV-]:+^Og4:
8>QY&<C,93O#G\.B/PS@_(b46/-P2deH[Kc9SbS^K[?HTGI0A.Wa+YQWYg#Ba0aM
U(cGFU=a[)]N8_F[P#2=4FMLI-0#<23C>+2I3E4RUO:SY+G]I95=1cI(FQO]<-b#
dEdOM&e;Y.6RWG@9_5+[MPf6>G>^@;MAQd&<],QeeCc-TP;48/F^\7Sc3MgU.AUK
4,;-.GZ+(L[[OX1P3#e)YA,70AYKM]EQM&-1^R^08]6L8Q[VA@^=7,DNG.>LN8#H
:L^3bgK=5+7#;,;E.&<PYZ_;=f6D[YEKJ^TbZQ0=:W;IIcf#;ZM[3;5D8F5M?c&)
5)BVIR1GPG[C8F/1D17>ONU^[JS->V2YJRd>&aLTS=aHT7W_#P_R.0WF:=FLJ_Y5
7UXO-TI,(6.gg+9g-a(?K\c#a@:BC6Q1;1MB\:@&>0DXd[]0+N\@JZ0H(B^Q8.Y?
8&=PG36UOa9(F2L2^JAP.T0TP0IIFcQ[bI#9LPC@b.AO^g&CG]>.NOTF@f.<5DTP
UT6&/]dK3cP<#C6FQYb7U(FHQ1XM#5XWcY]Q^<^7\d,Ic8[K/;A;2-,Ua4<VUbTU
2JG-/IS_(?7H),Ya\?_RBW&M,Q:)<8QAc6?DObXaXCJ3d<cY?Xa^R4>b([9d?6,T
5R>J-c;aR-A+UIgMTf^Ta[9P6=[R8aeEd),YYXZ0B17=^2@L=>W/ZH+6Y?_5[R5C
/0>S,b@@DE(S,JfVNWf@?Z5#=_=OFe+WN9eO3AR6#dW?Za/JE/J@+HeYb26UVKb]
RF;;[RK-fX5.^64e_B2e\YY.>TN8,4KL:8cZ\dU_Z+H03=Bc[GJDF.__70FFEc^+
I::]#]f[CQTDY6^&Dc+4JL?EP3&/dQdC4HEZSbY>GW,3]]N3W&9H>dKdV0[7(MFI
PK3Fb[1NW-a5DY6U(?Dbe)6YJ&XV&D@SB#NbXeI[3.FV(^3;TZZJ\^Ee2RQUW]Re
/.UA<FcMAO\7eVE:W<[RcM<((aAU8gF)RO?FaO/=JRN<P:d.1RQ;]G,a:19&Zg.A
..?e\LV+>1Ig_Y0f4F-XG=/LCbOAE187(9+gP+83KB@P<G@,[&YCPGeE,U,-8_ZJ
YCK.\1@XG]JOa5+Cg03<H7Z:Z(O/7MK9-S.@CW/e)60NH5AZc39<Fe3G.8CfY?V9
C);C.=A2Q2T-PMJ(@ef)\#[b5,G<Z+P;X@]7OeK>@9IR3fGXZ&:b_ZORHV@BW?1[
dMbd3V,-Z>PO9VeHE>aSL]f7fNXA).ScIdF[GScZ1fRS]e_E7S5CdcNe7?VD5JA<
9=M&I;JW(66BH7Y.&5Ee4<8NK(&.NWacbTRT;b#Df_L#M+OZ@cB0_VcK/\;.C>XG
=#KF-C=NG#VUS@[R/.I#AOU.)7dE#P-a2=.0f&CF[6-82YOWOgUc8#)Eb_+20\HG
)4JA42=Dg+HbT.3DY(WC)UQ<6A.@O.6eK=aR?[dI&:PMM06+Q]-dZ+8R?NIK0CH^
RJ/2;bd(c(Oe;@[PW)T8ZeC[ZeXeBcL>e8I3J[Je1]@(^We4R-,F.-Fe1Q4KBEXg
&IO9H@?b4\g/7^d)/FAVCQU2OQZIA/B>gMc8468#d=G,0@b6J@M0Pb3\,)BZ21YR
2/C<BegUY;8/38KU&4dQ>WRWQ/aM>YQ9?<FBNI4Q^_1_Ba(AGbWC,X9/08UP,c/J
O,/:EWBQYSTP#3_:3Z?U?Te+HI0ac:H)Y\>OTPDORI,7ffC/OeS?KL#f<;,]]M+6
<YbGfUZNWcJ(HdYgS\b09VY(K1PKLN&FH,&f,7<OI/2U.=(IH]d?](R9ORD\FOZF
_>S2_R##;RL_02L>5DY+)G5g(FW/P^EK0NKP9W.@8a@DP_W;d1V7PT2EIE^+@f/_
Y);6V\MUZ_9SF_9fROFXKW:f:#f(e01IJE#P9;&I&QA&4=B,L(DP.#+N;e_S@?V;
R;[V\>#9#d;(T+GKMM9\QM\5\,6#J;\H&GfU@bdeHJ=G/bTCY3cRHG=XcJC7Z\AB
#g/1[#8b++/IB\6JTeN72bM?E_(:@6:N#C.Da\-T:XeD4EN4U<cN[GL3)d)WI;8&
,Y^9Bf,d5aKP]N93Q</7d930A&[V+=fHBV_9W=#cG6-;GBQL>gGbP/?F<&cS0Y\.
Xe9P5U:<6P>)M3f:;aU1Ef,Y?8N0gDW=af;&DK7AT]5D)6#/+-6FXMa3XMdRI.JA
BeG<a8(81a^@4DK]OSWf[UQXIa=RFTP:4\A#fQ]Cf.-c/g]>UK\g,dK7gc-4bfMH
cWGCf_eE31>CO(.OY6/OGYSGdSAQWCR_FW87E-OLePY,8e[-Lf)JeN>=dXdLL5bL
@(K@1aRg/@]1aQ/a6Kcf.Vd5/,S:@S(BH5b_8G<@ECB1<UY#=,_WSO2/e]DZJJYS
:J[5,,(JF0N5.)RT:?F<+##IK(MHV0[=g(A\U7K[;)ggG:[.D_7-ET-SWE1Aa/I;
_V2FV,2,Q3d@aTI3++3&[,g1([\EdVKRGB9;?3;OUDZfQP-Tfa<U_.-KH,8,WVM_
0DF+/#]3[d6Ce:W>d98L7e0:FRDY+VEO9XfdXA4bO2L_eC#[B&9P;]>RIf,<-2c3
\Xe+@-5]IX/c6fCB#.02M?bd\db+7EI1d^=9CZGFeeDc/\c3/-;#\W0TA-(5R99D
H93Ta=eJc\g9dUK]Q/dg+X)7gOc]a2=92.F3d#TPXWU:JB9:/d95R<5T7/fgWMI(
XXIUaK[DQ.1JJgfN_5Q,-Q^bQKY((.<TPcMfAQKGf0\aE]g/2OIWG,=.G6ZH7geH
UA_H338UAJ4&Ub:#OA>4D>0R<aXLM(g?gf?^Z@:fNT1:;QUc)d<OZ\+H;L5D3dJS
=/PaR.<4S:P;A^4e9#G9EAHRKGAcbAf2FRH68fe^YPH+=+02@OKPUbgU^022P:N5
EVJYb]5EA][B#Hf58YEE9L9M)F]_XIe@&Y>1IBM+<#[\;@8+[=E1[NT&Z;=V?)/O
b&E_[7&8_Q2[2Fe)0G/H3YX]YCfc+FRCEFR[PZHZ396[.W@.EG#&:HF/K:OE^S-M
@TG:.cIXb?SC]=V[>dUU?Aff#JV(4EJU3cf]\)63Y[g44AT9)g--&5<C2E4T?WAU
=F(&G#9BC>Y=G907a7+C1Y+#aC6)5R?M.,Z1S+a5]D@aW@_:XT/BE52E[=]]CQcd
g.cMCSGf_C//EGW[Fd<LGdW&IQPBeCPf[\F7W3937B.,DSPNGC1;Jc-.3<GVG?IW
D7#Md20W@Vf-C@aSXIdE;Qg7Y0<3)Dc8Bb>LL[6=ZGgKJE3PS?&,BM75-]7S5cON
_8,@a67>I>WebAY\R()F#DUDU&K<@>IQe\[]@BAa(J3<F)\Hd6HA,P0J0Q&3?TUE
WITVZ^=;IZEUZ[3^B/T#NQ@5e/KQ)[Id.LN0\)_&5P^G[5dJ0:#R9-PG0>IA003;
.E@3U^>2+aZaJX.@a>g=?UZWFa9d2S<YQL+dV>Bg0\V51-XWb8_)cE(A\afa.X[]
\8WZ<gNRSd[b4F.NXOI&]/GcD/#5#E7.0.6@HY&/(&2?fU7cPHRXJH_aSI-K,FeZ
/[7/=W_(cYgXf#H7GROD-[QZEV)T(XBR>Ga>62N>Qd;X/a:g]LCJJ5>3&NLEW)RK
3Q-:#0/K+\-9a,;.I@LO[T/bZTP7?&3YQU5<6K<Q[f9-P96S\cNZ0WAGEDHXSZ/U
2^#S8-ZW062A<Q=5[PR1,H1;]6WUL(HZX>PR.P)b<0I1YdaRf(WQg53VK,RH((O&
+/1g53A>K(NXA)DJF59()g&\V>FS;T?&#1\Y-H:/D:BUA9L\@<=L^R\?Q@A^^+bG
Q8KENE#c5A,AM.G[Q+@gXDL#S6RPR&M@W=4(^[G62#CD.K&eI>-5;@5/ZC9KPU6P
fU6B/CQ&4N>e\3>?bUOOWTA(cHY#IXVY?Qg+=[BBM^@K_D@CVDGK:/Pg1ZgWGM[A
;Tb=.CHQdD4>75<J(C:21Sd.C>dT^bNOWQ&Q+MOWd#eHG(Gd,=Da/I:CgLcg/GX+
0dfO\(5(_:f^ZeLdI_X\BS#RIU07IW?.HBH<7]<_.cFHcE?^0:[K9,E^R6]4LF#;
7I/;fV<C+5-F4NH;</VX^dULDKMHA3LI2fY_GE1],5U10+UH.T7N@a6HX2T5033^
,G0Z&[AT6/^II];d@EM6G5SRKG4Hf1TKW4LR(@DJ&_#KgG-<CZSEg:.1A?2ZdB(+
>A[QA,KKBQ,);Q,&^A1[<&(?ES==UX^;QY.0QTTBVW3^W1<#f(4cJAN9Z6-<H0bE
R)-H9)/NEE)PJR@O;M1W>cW+P)_RZX1L-;K8Xcgc8&X00RL]1_W=I5PEf;5>H(;&
FbB9J4P5OXYB=-Be/R]^YCOQ/N<C6O>,15EF;?4_@;+7_>2^O\GO0^LSW/6/JFe3
)f_gLB)/bIE],5BdTKKgL_M46CG\VbK<@9Y3a@WF/AK_4OGPOFVeUK=.]/g5)d_Y
E.d8QYV,d4?XBNA5X3)5DcIKK87SW;?B2MBf031A3c1D/JK=OV<4:(,<0N-6M7f/
:POd(QJR,-P2f;\])#\@5FE0cY[f(5=SGT)G8NHQL&8fd,#AOaeM/RKTJC;9])g-
8NLK&8&#dJ+f6FL3,-57J=,a^@_MO1:?KMC86+dDPYc/bbR;V.a\)c1.<_VI.,2-
+S[[;BX8\:Y-<=&+BQEMUfYaMJI[-)SeO>Y8]E-YbXS;6SH/7-(KC5V8NbaN]RbM
,FI0?R_2WM:O[_ec93C2KXO&,Fd3gBIW)ZYOBW+(5=L_>TKdL[ON105_B2DMQ<0U
2XNf8O4A_R(Ng32M/f5:2,\dP7ZH8Pg4gZ9,S&0ATILZ]ZU;VXR&=a.0Q]FfBDW(
THX,O+N==9#DSN&)6.=T@JRME5,]BV,URaD.8S]_);=/LH0eZa?9cGH\[DSW/cAM
>I;:RHTff6SbMQ\=(X0[.JK=9=Z&?U1eX4YP@g9U.YBLHfHWNB2a\]J/;H])-B@]
=\(AC-/]Q-Ie^012RM8PE0acXD:HV9G=<2<RU/gFUL]U;M+Na<.&@LVQD_[0:/e&
);GS8Ee+fT4XI#g659dS@Z30S:M,bMKVSUE:5<N70a_Y^:#c@RMYe07Z51(9+5If
gPe++(B5F_RI/W0HW,;I]EOG2CM^2U17K4.ad<NT=@\C;8[4<A-J?L(2RUF,]8SB
bBUBb>LaH3-#CG9f750J+G3fbbfe+Q1gD3cR/I=#Eg-V7;aGd-.>#)QE=PeO>HY+
KdP<.Y3@)_\Nb(CJFP87\/4BZ<5I-&GVfdO3c[M]>OOKE<G5FJKd#>M?WB@&NP.[
@9QM<d3+(LeI?IZ;&=a,?B0T.ZG:E#P\_4V#LD9Z\85)@AP,.S61BI7e;7eE_#+.
I4(D,,Kc;.dfL^J0eC@bE/bM#BZX[AN>>OV2^[NSeDH6]cEB^XDP#H6PfVO<8C-;
-T=U4SV^LRd]N>3V7[I&+,S>[54f6;UR?QK2[RH#U3dOE2YE?WT/Y:>GEOe97U)U
@B)(^-+)Y.H>V/6^O;8aS\Z1Q],S]?YLF9J<(9_/I0)E.XOY2,8/=I,GUGAPK2cH
M_e#//e.=NB+E63/g^Ab9:H[A)8JB[\gUYR&0L?G4)9NAFSSGXL@UE&X=MUGJ/WJ
ET2K<dQ#OBJ4UX(T4-U91,]8Q>^&I-P0UGKQDHYUUdW@5TaY0;Ie>TRB:94\7FI=
K<Bfc8H50.72VKF?O2S],UM+HM0U/6A]aKM95W-dfC)SQZ>:O&:c/80E^.:+g.[/
N-:cV?)PBH_MEJB4;UF?IC]B)dUX-\F3G^O-cbGR8_@RXJ0A^Z-dNJCOYbP(W\?[
:W]J3b41c8HG^9d>W?FfE&c_U?.^cK=3[G/I>R]G+1f)9PF;/T<01=RB5OdQO1B;
XLHPMJGg5>#J?#Y,]e0#fQ5,H.TLQJ\(=PLH[D+8[gRe1JO6d#D<+SL.H=^EN+B@
+M8,;\A?+IX]+98P@dULNGXP6]=ZceKd2S5O0=ANRcYf\:NI9+\aW-SUg.H4\[f;
bP1f?R@>P=Rd//N7bIWG0Bg4/G1/<MI31.M@RD6<f40C?77W9CQLU4a[Y7\&D+;S
N>04D>1EcQJO/;KT0J>#&\g<RXMK?[/N(Ka+<J/AfAdSFVU8<MRTF@PSOIIfH.=F
=3G3O,>0&W?<eQ.^bB^YMIWTgV?RM+KL8GS,dAJF0#Z29@-DE1UNX;WZ,de7G(>V
3/([835f<:0V=5TD8\b5R-GbbF&(_].QD-_dUMQJ,fDVJW6E#@Z:3>MY6=0AM]ZJ
D5&VC[,6RTId4N]@G+KOROZ;+Yf/c7)&Z\9;<W>#^KOSLKcaL[Q69S,c-Tcc+[UW
e8#0ZIH.O>e-dgKJ];U@#7/G&)+XIdA6<LgP;DS^0dVN?DaEDRF9VMRDU]1#C2QK
0A=X4g-BSGFZ2Re(QE,5T:\&OdbN_gK,;7A\6fB@&5DY?@X@BaN0(TZD#&7D1IE#
JL^Qg;:D6\ee8Q3XP4SaW(+@KbGV)dcL26eYH+_?VV9f\^?<JePJ<MTJRcF4MWI5
0HJ3OST#K99301\X-XY]?a[V;AIQ,WQN[(RaWGdK/eVUSZg_^0NFY&TQW3FeK_.@
;J5U.RY95Ac6=&VCA8.SW=YBPZ_5FXd\_#GRVFD2#bJUA6(Ia;79_NfNOTOeD.+8
=a[3#EVVP<NHgd:S?Y,dKTK&bOF?-(:NT@TGJY3X&FT7\+G9-V-VKIdOE<S\bLcf
XDV^g?)6_@^TU5<YZ[@2(?3=d/T(AQBEVL^DRbU,CLMH@?R1cM4:Z&-35\WdR7Za
>bHBX0FLEV[K80@:e3H93AQZ&Q4S3>[,+Sb=C6?OH\OfI<W>N&#OeV^=8+#LaT(b
/D4DPHTIaPd.(fEL;-(6<Lga;G;?QdJ3RRWBA?&2/-\SGBc3B?&(2d9gU6,H@WKd
]W;952g6S#HP71;YKVI&_g4_WZ[LT=#F.(LHXO_+)bIO[#5AM#;[gQb<T9\d_E5N
X+I^777Q4_7HWQS;KP8T=MFREL38Jdg1>=?,;?cX/D4X\5[<41P.1.Y=?7Ta?@4a
d[@E+H?_QB;J/,LP7X=f(=d/G8W)R(9L8c^IXK@_&YEE]52)J=^0RXX->b#_9VHA
>LBaa_]]CW)KUaZ8g.e@L).@T56^_+J>8D7->D/,2aMbRPB6f5=><E-2U1b]^(G/
9WdF,Ya8ACE;2R;D]<3AFW>\S&=#9c_(-ED.FBeA+DEAJTVY^U]f5V]U^B,+B/I1
))_<f2M]LGD&BV_2^NaOARKSLf>:GER8W=UFK2G2NT^LZL:+5P&)?\8Qb)fGNTF/
HF-S#T=\F>g=(J01MT5LS3d0E?1_G2=cN<a>L^fS(?_d?R3b=727;OJFge^5fEOF
[D#APV.6MBaFSZ<Hd\#]^aWHOA^fP#Z9)b?/eb>@?c(MYCOBU+==[^;B21@QF;)H
YT:I88BCGc)Db#6L&S#Zb5R/7E6IcWL5EX0a_YNcZ?/EA)S,8]3R>HKGC]SdZFC9
57\F0/Q[U49),6T<]0(QWB84.FT-7C-\>f9JO9cQW23H?BA,e:2Z]J,abD:9[8^W
Bd?ZOKR<c-]FJZN[fU=_4F/cK=HGZF8agPGYV6Wb+<&YU?V5GS83XP[Z5;B@@L(4
bR5)DEQA2)QK/5E;XA,cYD<AT90UB(Q6E635PEA0:&]TP(1OZGDe1&fX7H6Q8YH5
0^A.>O<=0OcPMc=B?R@KE7M0b_CNIIeK:bWEYF;Z=NeY-c.53/dN67=Gc?)Z9^.+
_M4UF=T]UD6_J4Z3eMZPA\4Va92+6WfaVI>(9\?.3Z);ARb(7[Z=(BYM\L5KB4YX
gY1BdUVJPdIR5(A?#X0VD=MU=7=)&8BBTMZY87GY>X^W-?G;CXZX)?TZOKc4VG):
1IF0L4&d=8^_)a>B4gM.QgA6WF#D>.S)<?][=+U^5NIZf3P._1=0,YELYBf&1B6:
LcGVY[NYTI64E_[FWJL,OadWZX(2UAJ3OQ)T2CNNP7/b#R_GDG+/2+>>GZF<bf&<
fNA=Qb(^6=C(9L=<Z&f#7#c:T,4NSKYT:T,-J:Q[d>X_VaeK:J)J^^Ig0.STYQdU
PCZ:]((\7EYDeIQ&5CB8XY#4?(THVL=BJbbB&/I&Ea1gcY)SKD#>?]FPe6M1S5.W
^5)OIE?3cTbEKEd76\Ff9A_.+AFT@<]BB9Uf][)BFT\DK8gJMY-EK.CS&H:6=^_I
4C)42NOLDMgZ:,\O=NYYDdEZ5398+5cXKO[#I^^73QU<X->Ne0aCVWH-Z].3g-=F
HGJ;.?CX:YbBQUQ+=ONb;fO_WPS=PN-O>[A#CHa=ZNb3WEd[.HMA.AcU1P]FB,]d
99=PF+S[VYU88Fb4B5c&?.SO<0eM-=+/cXaYb>/U/_])(ITKc=P(/^J.Nga7H&+G
MbG/9_CGA>3S&5a[65AdL:GLI05fDVFY6[I?T+@-aW/6<H>B^5^5MGNQL-&[baG6
db_9B3Le[E#OcG@\^RM@WPW2+=_6JVN]H)FgBFG4]?KMHIeT[He#/[1+GG,[BSGF
Zcg(C@c0D\BQ,1WB+7GcT#_(7G#.BHa@-+=3H2>)Z=7U9[(<[VMKJ33R@1Z@)5Fc
X,;Q)#fDf)&JR^,b^T3UgNAIM\VD=6.dG[#=H&J.PKXP;G0I#+eC:]A?G4d9.VXO
Q8MG9C]d=(Rc@\B&0=S&A0><MCa+3DG7>5WF017T#O_I,19&6+6[QLabG1FgHBX:
<KB+TPR0b)3;3E]F<#;7T>ERgZ\Y/NHT_?#B(U+&:4]-Z^<2ZfHYP&-7S=A?9AI@
X-5d;/OdNZOaY7NG,QNf;ISN:WU;2-g6aX8349YTE\_EA<gI<JLH#WaMWa4S0_C;
9JC)F&MgfOR7ge-J<]46@N?&IM4A7gbeM(<I5JVa9a\XG6>.L_,;D1XLN65=Rg_3
OBK28W2P3YVL_[U+SMJ)<aKLL)J#_F]ZL<Z)J;.c^Z;W:Q^.7/FccG?PZ=7?H>W/
R(@03NB+A]5D9Tg@6Yg-YB3R)5deC@,S;&0cLBWSZW?E&U+eBLde=e,WST(O>D(7
Hf<,^<c;U:ReTL;[QOcc@ENa0XBXC3N,SaO+a5Y,+JaAE3XX&aYG)M;@E]SQUXD5
YX<P\XJ@(L,g0Keg?ZL?a>-]U:cVEC^2PM(TgI[cQ:T(#I[__CF:]D@3]KMEA4\g
3fGdNX26?IZ\G@b_SJKL1IKfeMeDO,P(8Tc=IZ@g?Ag3E?F,H&&;?Wb+0+76G.GJ
I/_fB(ZdVdefB.A#TL:KE8eV_[9<8R[;.9.0MQS+Q.K1@S:-_D@P_^:_2;R1P;;=
[7PM6SK[aPIW_:F2T,Ha1e9@BE]^,-(46.P8SW(KbF;G?\Sg.4?1/Dc-&bZ6X-L9
=\0+[+cGGW>;5Y]f0-K7[_UNWAeY(-;&#PBe+(L38E<R+8DH^W,<aN.bdT6b&,NB
C.<G^[K.SKZC1>#(X9:B>AMC(CFgHe]KQL>XY^DUH^Gd\T5P8C50ZYJ9&+NVdAQ;
X6Q7W4cFQ3._9^B0IRc;N7+;N^E:<ZX5L,TD@)V3MU:?/\]5OP5N6..IC47:2XZR
,V):4[O3\#78W0P>_[g.E]LQUAdB)OM\#F,edOX>^?DRIDW+;:&2NX0MXQ?g)&E)
VbUe#Mec3Ud^ZB;acIDN,7L-/>V;UCH&9HX95@?K86LQ#9A3@9HWDF1R^X8X43=,
R-:?6=M#JSCIO;BDFO&Q@K??#EK07&2SK18RVK-Md2B5-LCA,3dWb[Q.>Reg/[MH
HM(>ZU_[(JD+f82&&)G>(408]0=I6EfEG&gIZa=2;VBQJ1:B]LO&Fe8PgO)e4#&V
U4[_NdY2gQ9a)_RBSeS^JL:C3.=F/J5cSX9:IQZZ[I@V=>DD9KAI:9:/#cAgGT@U
]19,FI._N=)M??:P0FSdOE6]D1_T&-Y\.\B3AF8._Q>/0:>LM(JGI28(RV#b_eU6
gKD5Ba,KFY0J0]KLRe<>R>AWcF+#GY:@GQH6;1Q@P#ZJ<=J(1XAUT440d[PbXdP,
#56BB3V_&)\P,.9ZdRa1=[>L?3f?dRA:/-CD0HN=QbZe(X0I3[-Q]Wf)e6GEU.W<
=SI@GU[GXFGQaA5Q2SZ8eH/>@K-JNU[JS@f7-2.AC7e96RdL)^./#YQ&.;c@09\c
VC;OdV-4#;Ye,4D?;Of0L.RgIK,\?@WB9RfX&a=5=d)5bLMIE3O2>HgJ&SX?/_/0
;dY^IDR6S>gA3(7AB(-X[NX4+Q2YA)DWGdMZC@9FHI93Q9+4g_EA(RV,H(ICDa8F
9]^)#4f[3NUB@>I5]:(Qd3E]=Z(;JSRE?e><FN3UT5;d^fb3DLENTH=5X.W^E.6@
7(>IFQ[+<^H/7/D@]Y3/LAAQ&ZK@;(])2MQ,O1EfL1UZgA8PB&ZJa_BP4g<W^.cC
X6<H5TTM,7Q=&I_>8bIQ4=:KdWVENDIVVQ#G+]S=9U/f&?3Q<+&5SU9[c55A6A^Q
TEeY?QbIW-3=^7CFfMSH1L95G?8;gRNPM<7Eg=U@CPR\a.MA8\Xa>(<RAG[S=32>
R@Q\JM(<DV2XZE@I=<LeLK,[P(5PB\FP].b0g[2VO\eOU#OOK:f3#gUCO6J_YS3F
_,b(6<M,Kc4@?U#R1>BUH4>Q0TL@(f&WGZ&?-Ia289;E\Y6fB-FMX-XUVg^MHNEF
(T.YaY)6GRW-OO2^CR6BK-E3K>e.WXb](WR3Te8E:cT<F)IN:f<K#-6ZZS3HN?L5
,aScdXACdc3S/MM#YbT9/[b&/RPBPaFBd)SOJCB+BI:XbWA\UTON^IgV&(=0DA]N
B<TX00eb\5RLf7832.c076JY)RUa^+SKG9JBM89D#T.[gDJf>&UMb]U_I;UU64@(
:W00]S7Y(e^V4)1?SQC)g;#Kb3b1E=G9<D1BC&4eNI]O>7I#?4VQ-g6:V\80RRSJ
eNDdF1dd[9,g[@RI3LTI^7[P9B:5X]P,?SXLA;egL+55Fd/CS-=-f#R:[e_],=,3
SP)/ACG8ffX@U>JO80IfS3I>LCBd\L)@JRNW^YgVBNfEVRF0Kc@Q9L:>\0d;gL7U
,42B:=Tg1N8^GXObL4?M.<#LZ:)gF2@KKLN5+CQ<Df9g6IBYOPYW5>Y\2OLf>/T#
\YQV\gEN++6fc5#7+<RY(+]Hf(8@M.KGRR,X0OW[ER&(C<\8I?=Z4?KBWR9U.7ZZ
H3KBCM@@8[c,7P8AQ7:a7T>fP76S]5#W]4[&5D4>F2N\cH]^(-:1_e.4P6+KV7)+
EB<@-+(MFXg5Z3]T(^JQYX87PE#6@XW2T-BgbSN9g0SDJH9Z?,gY,5JO[+d)JBd.
bGcEZP2)0^dO/;]b1]L;e:P,Y330JbZ=92\GL@:_?=9HPB[bRG3;aA[\7/c#@\:J
Jd7)IfO)+)(LS8XD[EY0,)5CJQM;]\2AXg\_+^9HdOX:ecF0/N:2,2;S33+^cUg7
g/E:M?[</e[O-NHT10_JBfK]gc8N6A?L1RYB<?SB,:0\[J71ORV()7I&GL;[S()V
LOU\C+g^9#9KCTUQKWdHNA:DP)N[#R_;EY7X0,XD#2X/N=^8eJ\fG+PKg\0>>)RD
<;SgZ[>,]M5Wf_bZN,Ob4QZU6RC<,I=8e,O7-V;7-B=EGf^bSWc7JG4ZPGO,EI9;
@g7^7YedFC?VV4VZ8./0?_e)gH45KZ(f#KBRY5X>dAC\?<YaD^IAEPE-C#f+fHc4
JZD0,IcU/HMGFB>7]V,372:^BTV+0M/-LW0Hc.HG[YGH62YY[JNW9V3636AUe/=Y
3)Z@0T3S38FHH+JT+/IT?7&,TX0gDBM-)CGgV?7AW_+G5=6+V/HTdG8a+37A,<YI
Q#]b<C0CXGa>9\\FJ306UY5QF+[HKWB-,Fd5)WL-3ORZ9380VX0/U+MANU2dcXD[
3Eg42G1NA@S)]4HJ4[2,:O#NV6I-=J<]8=D-8;7O[RSC.=/H.F3^@&b0(aP0FXT+
IJ5KD=@A])<5?>/NK1W<A(+d-0cQ#.#>TUOVT.MWKFdLI\DO4eI-G;4#](8?PPUH
Q,(R>1[,=R16VO?<U7eFIGHA0>:;^?7C@;X/H;UJ2OPXCdVdL]^VQ?(DGCOHc3M=
45MA1=3NHb_P548B_+)H.:/@RI;-&MdA=#FL.81GGTMNQ[:&^2_AD4SH@M):\7^R
WYY4B7b#)A4:PP7X@K9S;eEA^f_+^BF5(S2QWI:D#T]=cN2FTbQ55Vg4faT.\M3,
HY\Pf;AVIg_&W3-gUV6F<N(AYB5/c]W=b[6Ud3^AS=K7b);Eb4:f/6]\J^JC9?F?
+,?IM/<H2F(MEdM>38F6_]MPB18YZdd=OHVND65B8QF2_YE/R,<:L29DM,@^YDD<
a3Y9M_e?BR/XH?7ac8[,4(XfW8D.KUQTLK8U(?KXI=NMEcNZUb(g\OW&0V&DI7.K
4a2cad4+;,YKQT:a);U(8=gZN[M(L-W=4P;QL)IE@GIH>>RA:GfM^fL3._&WN<SQ
>[C>,CH9Lf_+8]L9gY[cP6@NH8TS;KBL\6?Q[bS8S-Tcg521ZT;aW7QCF&U<E8C)
Ya_Y49d,]gM,0[+FQ(DbW_M4JTf-dQd\@:R:PF^(cg[YV50M/a.XF3W_W_XJfDR&
H6^7[9G\T2;Y#?B_@[VJ>;bc.MIOML.Hfd[3=E:?PA<XVd3a&c(UYV_G9?e[Eg.2
1K8<F8>I@2+]M_MN#P@G(-3Y&L0UPKQ=e84;_Hc&UOA>F_.G,gY)D8e7E/+ZdA]3
L_/Y<TQUI:R,9:)HI99/.C?DeA56^8A7Y[^=^MT+-+0<KSO0E?IC5fd#HSER:Z_f
UAcAN:d.c?,:CO/#MTaJb24?#8d3E2><E0]-GL:FcM6/f,Ta(,ZSB]]f,BM,7B8T
.]8^fG16U&_feTUg]OZbP9K1G=a\&8HS15-[U-9C)H+OA[)P+QL.FUFABcTg5T)G
T\:XC;&Z7IQ>-0(M5,9NZKI@-2^H5I,?)DF/VZIdSe?cff_>?Y6IIUC?ZQ9W>T@(
_HaeWdU8aXXJHOBU,8f@c(c<:R-9PU8F[bDg@S4KE&;FR,)9H:1bEd=4Z/C\(9&E
4Y792Q00NKfW9:5[=T\GNA4G4[XFgUI(0MDQ=@Y15Z#+EYH);KW.d32A-4@AF[FB
5S:9e<B<)U[6\HGIgefbGV:d#YFFI.K4DY3G^9&#DI1AA9N:BMQH:A7#[IM+;1cO
7Bg\eBLAVa84Y0313-\7c40/.-F/E_3X,F=\6>[<0\6=c5&L^JM\a[/46V/1gD8;
/O0IKA5##><=\)Q5S&acFbJN/aLL;HS]_SHE(&V;,^06<Z2AU)GSYYMJCLcAb2G/
@B\D),bb,G/UH+Q>R5C&#9=E4RXC]+AR#&>b@fKI>..G3.+MVB^CcDd[&7?NSeP7
KQ<Y0B,#WSCQLaF.e?+g6?:^3UB-?A/29N(SS^N)Y@CSPQ3C6N;@^PZ?ec=S>bDU
:K9KQ\?C?SFF:34Ae<-WP_?ZUfSb&H)(SBG+ZN0?P=/<?^NAQ8]U@d>;#HWC96U)
BF9T@7f_-TegHBCXK@S^?F=4I8E^;41)IGE+_9Cg.\HGRT]5D#=,.JTS\6^)T@M_
P6M>B,53GBIe&HM,]&.>e3BG#@CdK4/#Ca]+B+^:.>(D>/5(-e6VbIO5(;O@P[FN
f3.ZQ6.>_RGZP39b\e9a+bP[?JLcgULQGYR_)d#+SaHa2:VDGEWIXJ_W:[8^RG7X
4ICY]X:/aU@UB2JXdZ8/bN&-M#:+E3eSUbFJ0IDa.5GSUC:S?>RE32gBf5QfW+-_
FdA<KDN58dX\Z]-I#f4<2MM?CT#6NSK:Me0ARAYGNXK6[cYLISd<_9e-8M[Hc8YT
-&Z=&#>+I::8O\:Oe:\Ld>7PAf+X^ZZT#>A&_&ff2U;;ZQ4BW#XFU;E+(1WfPCF1
<c<g/KMaKd?)(VSb8fA>2f:G1IB[VVDG6EMTCQ#E,LM.@g#Q@9P]\@bMV\0Wg#R=
/88&<Rd^/fJDGb9WTP&]1RNGECY^-cB&35G2WYa@dIXc)H>)^6J;7LBC/e+B=3U2
@)DUIBa1E@eTAD[R>P1+d<SO7B1bC;d<[Jfc:9_]UR\?gVP?_4R)KQ.]WSFJ,4&f
8e_5Tg6D\R+1c@UXdP,(_cT4]87d7=HUKOI?8KZ.+8ca4^3OD(HL.O_+W.2OU:0W
bK(7:1-XV#,4A#,939O[abgY@?Ceb?:</<=/0S>\_G:?RVBW+\]?V.T0C[YC]#bT
E3)ZdbFgSeW/Ad[.,41,A-;F/Y;f.IG>[^b+XF)@S[WDA8@>XGIKAaZC^c)L1_e9
ITNaV?,[:]/,gP+Rg)[)d.U@T83J(BO89FR__/KH8<^]24eVf]F>>\C>N4B-Y1@B
-[=>gM/],6X-T(3>?2^Ta84,RM;9+&70,.LLLUJ8:Y)^SMS;C3R8^4<-79fWEgO)
B8ddIXH(I9;U0Pc4UMG2K6F>0/PX9+[;;Y=00-\YSBV7^W^QgU\a^7bc;_6L[Y0[
Og;0:b;;RNGR<N((1_:^-(\?[60<XT[@2aC24M-=7=Z(AP&#BC?FJLC1Z=P]fPI(
@I]7R,.Q&<)GSBEMI-\H336#S^[ACf4[VUK5?,\@@7gd&#e\B<CK]^L6=+]IecFA
gCMZQIgc?D[=5;aggXB+?W_1.AW-CK1_#NV9^\=SVd2/-e22][Z33UEA2S(WUaNQ
&1]LHUe(J.0G9_1Ff^8E+[J\Y^4=Q[R58YCXdIU@ePXRM+WS4c9S2PV.G9/4Le-D
(770/Z>Z+G_N#gYLDB-Q5cfbaRG2Kac/)WBOHA.g/>d4K^QMLf=c4T8ga7(^W]M-
E54a;QH-P=5,?IF:fGFI-URK4d1@;A5<7c+48M:8PUd7^C/7fOO?^F#SY78_W(e6
Y+\OgPd/,NV8YPWDK,=ZF?b,EA9M-2FBTV0aS>_0I)a@baDc=?_M-HGW\4>1e\/;
JF(8X3X)/5=[SB<a?3CT2KVSDD5:4)TbA<-]/:Z1L#W:fN76PWK:X\Hb4@JZf>HN
1MYBTC2>EFXN=1B,7L6N@://LLWWd7RN1H(OHL:DA(.d0A\X2Jae<PL;c@(_X23K
WLK6_UG\^OUHZXOFB])ZP1U-@6VG1?=5QeB5IOLE3R/TL3X>C8@a68E;R(Gb8gO@
_F]4>[\=aa(,2_c3QXO,DDag&gKAEK_U3XY&?aIKF@Af55K:b:+aG.#Z(f[T=@2M
WK0b0[(g8,g[eCFG[3B]\B]a#](]\@QQ(=5<\X\Y/1[M<.O7#6=8V=VL2-Y1S9aU
@^+M(R,cAH:@K<YYWPXPS=6M=PP^EEVg2(JAQd][;F>H.H3a=WFQT/F9BBUET<Qa
7M;LG[3.T#[6S#/05NZ7[f@3^b0(98g^>&_BcFVQWO.3LH(W4BK.BS/_R\)>9#bI
M+SE^1):Q=F:eEXe)RYFZ2(YQ@,:W>)f:,9&DOL8=c7N>Vc^3f.6VBQBP,O&ddLA
<9-NCLF(YdYPOL^M;R+@5(M.c)(fB;=]ZQR#@+U2BJ+VNC,C/c)HS/8=W2M#Z;E\
TRG8(baQA/c2Z[J2@ATZ,0Q1(T_XG2)RNK]_6U0KH)fU?f0,4_gPD3eCXK1dU5NS
&&(-)bYH>I,=FBY7@Q7^B=Mc:32Jf]0103aOL1cE(b;J+3DN?Ja>PXD[.R?f]1f&
RE5Y.Q,(6WB>HfgL0Q3MDAdJI62;3^YE9^^&--c/V7\)4;X;TD2aCO\aaBVYB;?b
_+BL,<&,W-#>dQ>R+Z^;,HL8SHS,M<PB5DIdgC.JLKU>.C^F]3gBX-+gE\/=)?6d
I8KN31aOG,<8HdBPDM#H=<VP?)-C+2IDUK5Y4D<D83/9\P#Z_<RWP#61VE?_JSSF
Fc6=L/PT-]KP>8@DJYQ<]2<SSbCNB+5WP#GegAWe&Ic;IK)J7F8BXE5(b1;dJ-/T
\N9&69Cb6[:O#Z40A?RfLKAX3]K+Q[GK1GJH+O?65:6]f0GO9I)@19UT+&2Oa/3F
2IgXZY[\&7)b1MFAAYS[A>VE676J8CI5,)\O0:YAQa4JXE0AWIS+4\b&,]+UMD?.
?)EZgBf@b?IB,O[CEc>9DQMZ#/P_.dg:=[?:E-HQS\;XKb&T.YR0.g=M5L51E@U^
.ZFU@AZKN.>I34L4^^gL]S^:2M=F773ANDNgVWc6CJ3Id7>(@E;WHW?\JF;7-+)@
(VF9S:0:BT+.]::aF1A^F[^LPY\S&[4B3+3eT)Z^XV:C?bAADG<b@E:3<XbF/B1^
L=3_3H0FFDNE<?7P5D7LXH5<fN^=TR^8gg2W,6db.=):f?JPWF(FRF>SEU?6+6FN
NTbPU6]4VO]K/M<8<[OEV\ZaJb2dPVZE.,e?0>^V6WK/T07\dU^IGZ_.W?=L8;64
7-RPF:(<Z+FUU_&g-7<Nd]O1W(GYEd)&P?bfa0^bB6V<S/7_MQZ-NWO#-f1:D^:F
&B>.5(G5<\1/Qa8fDA9UN^[T#6a^2(@?a\:X-[]JC4HRUS0X(d;WN<PW:a-ED^:e
VV,a;EQ^/DJ3GYI7#7\d[N5C4^78g-W=1,dIUbV#IM/\eDE4:GN-,T^\b3@KOfbU
bMX=OOGP5.>LQ47\NHK-XQe7cML,0#LN&+aU:#9,K:BC6c1Z,CcHJ+K62BUG>a]B
T&)D;2gW2FQg;bV&9R.98;e_C))X&.A\YJZS1--T6GNfAY/LgV#.+a+)=8#+;aK8
1=N5(3PbUN[V8c]5.@fW3NDY=P,d)^0gF_@@QeA8a<-R.I/YZe\GDX4,@MaB2B?#
><Dcf;YA\A2WZ.1FPV[_A0;(/DCX]NF0H?7IWTV^ODLWHGBM>,f]^WZ0<SE#c^gY
^.?HZUP8e<OYHOe,JAXag.(O_)T_,]I9^3B@\E-0F>=KFWVU;TJIbeN[WDeB7Ob+
g?9CE4BNMM<0Jf<2-b-W//d.&e41P>M,+7NaS6JCN-&4V.1PS\0cfEM&[W3R9;IP
a&/Wa:;,YB&4AZI<TYfIIOLdICa48>S)9/gQD)gN]8<K09>0de+^C0K/gM9;RPYO
#RTPSF[PdYX#9eDJ6JL1&cB/526E@([1;.a/?:7IIPUL,R[f,<_08Zb+:Z@^cT.#
/7Fd-^X:\dP3K80cVFJ;[<W[c8cZ=E&MUJYT25P=(bNH[K7+_QE_Xb5-=A]STZbc
PS6gY>0g.)&@P=51fN?gC=:1:\>^A(1G1;P#[:IcFd^B5EKd.KR+dd0bEPbg#JV[
WAT/?Q@U)(=g.?TbDabN)D1U56]KMfdN>Z6LO\VN&8FIU)_?X^.;ZNI4JT:Zd/@,
Q1>8\K5L24&,DZ7.7&625=WfJ0T81g\E35,:aUfFK[T.>C&4dYSXW]gDTV2L=DDB
UH98.AMD-fCJ-&.?,U;DXf+BY(KfD,>-M[::L._>U&[SgH;DPBW=&A9\)e];AJe2
.>R4A^?8F&0@PgJ57-=@PS??)bGVHV<ba?P+9DL?Z^P2182S0C9_/5BOCIL7VV1P
8d<N)&.FZ:@X&3)\FX#J+[GIgLZX\ZNM2])UB#A,a3D&5_;.570NY-N8ORT#Q76A
c1.1e\GSbRd-dDJcW7B=02NXS]g;QAT&NF3]/XP2F\-79#K,Ia@==KQ=<F<R9aUK
=EC70M,GIbR/;&A51Mc1fP2;H<F5.bFUG0A6,80QG,QT1M6@BTaZ<_:TPL=8]VcX
IS/@H=a;ed,5)Q@4>\N3B9193@e##P+LJ6\O0C+B0(=6cGQN6H&:AE5.JU_d<ULD
]57G<&1R?+7Q:NZc#a&dfE0EfbH,,2NZ4,L72+U<B)fO38@eeCZ#aLM-&CF?;YVY
K/)g#U+C,e(c21@RYLF/HX^Vb4W=R:RJ0AGO3D[f\/57\aedZcT^LWVI:>E&B4>S
1+S)6-&4:#^?6>W.?5D^SJ[@964<\b&86Q2VESD7.)Ba<?0.e1EH<^DT_Dd.b[fe
R[5JdF)VPV4;1RB5ALK>5e2;/JS&.(..A8KG[W0Acf^>>-Ye61Fb&J9e=J;\,5CW
B3eRLD,7]_T_eDR56S4a-)QC2H^K+F8dIL[cNG08_7YR2MZL.<X]IJEeEPa>@N?7
+=-?=^X>C\8OZcb>>5RWYC[<a.g>394XW8D_b,A5PUX3:0V[e=98JXW2E>ZQ-X]R
C3B&JN6(NM3a_,712CW.ZT<D8Rc-O]PU9@?>AV&>E&4?JD-(,:Y27<8G^CWT6/(=
__1g[TU?BE<-U#R>UR)=;?J&AR5H2PEF<gg2_J]OHcDV3X+YPRLL)0HODda,ZJ2-
\/f0HLd#(#D@He21YD7IRcSO9(//.@UIW>IabL_YKJ5WISUa/O>J,2=P1\B]_(K_
=..5eBbUI6CJTY[7B/AGgcDfY6^X.RNH2F.cI6HQ+XFDQ,W/5fIb3.LA</0B8Z?E
b.\>,.9IF.VRV@Q]gd.LeTaQ==93.Rg(WJ((CEX_J61YU+LXC^?M<O&;<O>,-Q+G
,L/eMOB#,dL9a8@8U+T&:4M2WY=7GT/2Z@[Y_^\2UK;0IN2JaUQ39RXId7C<UC+.
].?P^cD&5_@G<3\\H?f#5C/8E<_WJ=)0U2?/9L[I-2&bWaU4:S?b81/:,4[(31]<
Qb>M\2CO^3X[3-<ZgFS7N>V-^0W@#G4gY0b^)cYMAL6/dL9>C1W3ZH;1+K[S2_W:
OG0:H8O/(/4:)-;5W;:?+ARTZW(@-IUNDNQe6?fAbNdSZ]C[E07,bb<GK@[(&?De
bX9RT.KYFBFdg&?A[U1U17WBT(H)I<S2HT)D>cQ>^_FZdIWPA5?Z4\\V^6V-)Xf<
&K<a=A3:X2#bAM1#GI/4=8SeX9P/GHd7ZQP,[B&,S(cQ(Q>.1cUDCQGM@/9#(GGW
9K)fT1#U=UJ#<?T,MYa0#d@M5HM2VCJ<=?@d]>4.-Z?g)f1)WWg9/7XJ+VDH;5XV
XYLNZ8-0]0Wg@UY;eK1;;B>(/\e9XWgd.)f&PXD+g[0Ia+)EHS#&DYUX?/V;]Z<b
Ye,JWHCOg/R1<EGFSP+##P7YNC=BSZOWJ9OD1?(.f,;1-?BDGCN@U314__).C91R
7\S.a.9&RfG/IE6fA<XRRCPL[L^;caPKR4F^15_3G=))3R:Y4>RV6UJ:Q1+6b&?\
UO1gfcPgLC2MJe+^AMgc]_9R\Z\:R0-Te]E46SWK\U>?cg17W7f.E(Sb\_eJ8W<4
9>T/^CC4NGFQNW[VN]<J?>5P?d]L(C5NC<=GF-)W5,b4O5QNJ[&P0-^&;gK?LN@=
C^P?2H0_,-Y1@,W/eOX[(L-W&(X:YE7bA9C;<cUN6\K@CPEf9V4A[5W40(E\f#[E
7ag]BADRZ;)Jg_D<<^K#2PgOQ^@1HC.eUX31B8F:0MYg=GGdD:HB-O?&V7EYA.EU
KNa0JXWB=G(AF4c;bUa/&XONJ^^;a[[IOS\<AD0_QEZY^VN]BC5V\ZKQH)93@c)#
9^aRU^d&6]Y/_0dd,O3IBQe;JV3NTY<,8Bb>:b4+3F]65LK-E=0g)E;-[/YXbT>=
\geR/DL?AK.BK;f2BOC_I-L5a6.efUGL/J(P+9@R\N?^;G&49L9f6)38^^<I2Y>]
:eA(5TRXTDWU+X@B.M/=;I@EbM&@UYH@e[C(bGN@GcDO&QE/\(P4\&];C.;U6f1-
f@YE.a-c23]&BO^&9FOB&6&4O4:6T?8R^<93GZbAUY^=PD?FZMXR#12eE75+K?L)
70P=E=I[,VEMGW[?\X6XR]@f^aQ/(]/O;:I2\VUKX&<^D3K38/_2^ON,Y1e.cR27
fLG6f,A[K.IT:bVYA<[/J/[Z69WZ8.GR>N2P\&gSU_=97NKU-^?F^IEE14<0+gNb
.-=)d&E1;+8+Y^CM<gMK;R>@>6?[P3A:16Za;;8;PCT.SSSV4(OeZ2[WRJ>Y-Y?g
dV72F=).M\&9J:f&@W/W6#fA0K1b#0aY165Dc3H:N)\^;CV74E5ADXgH4OP;C.(I
<SN6<(+0bR.-ca)5fVKA4QgG+59P;29:a/M_fHZTfF6\gZOH#^@S3LDgGBR8\?c]
Ld2#LES2#ID7L>;NLR<2Q9:(.J342gaN2\a\deCX5:J3N:ICPP[61DN\L)TbeFAW
Ob>G7JM;IQ:@1<SVbg[8@4Z,gOK2N&IW\dfA+T<C&T+eV8c@N@9M;PaR()H1fWVQ
9c/>cPTHI>]3ZR??=&SFU<?W+Zeg-FK5;EV.def/aCO]HJgFf7P;,IgHIMQ\5&MB
ZB</6#K3]34R)\8@e/?=W+OCB-LVC;F&g9fd1R^Z=]0bP(8UOS-;]\b>(=DaHYE+
;3=#;S8+,GR,<_S)PG5P(CfI,RXgLLb-Y91J4>N[M]P3#SJT5BGL>PDEK0Tf5HF]
&K3[?/L;4+F?aXQVZK\^#H7(Lgd1^Y6IQG\f)5^(eXc07Id@FT1Z/R#SF1e@>KSR
Ic,.]_C0H<#QY.B<\QFV<<7/MJ3=Xe>6#\<U0cX>f7gZ0ZJEd+B0d190b65F?CP8
?Y-gD,S[24\50-\EMN7BN@B[>Q=79]aDP_<&]6FN(-US+>+(-(S[9Y?]<XPcIf]I
S&5LGBT:C:I4+^f,O6@]^F-eG<g.S(+X)COBT]97=Nc,cMC<M>5&K-1;#YA\9?#]
6g8c,[4fbUS0S3dVCG#T3[Y7CbH;&#W(K&65G9.a6I#^Hf>4F71R[[O24YK+V.LD
81C/F1?@A\)(GV3,&.3_<c.CQ/.(XXC#O)E<?gK^/<+e]\:V+fU>#4I_)1057X@e
I;H&?I,_CAdHPB[KA5N7L;LSERWX<A@\9M6AgJR)46G(?W9U7U^6FFAASH-,F\4L
JFcbMN0P[,79:;C2Z#H:0NTGJ,KSdgB<25((NSA[3VB0ISQXRZO?+#f:YZ79M5.:
B29g3A+K]XdG;G0:U<+?B[Yd;ec8/Y035.]+F9(Qc8R4?9Ad3O-2@[efeFaJ#S)1
CZOTcY?Ogf40\LV/M&(=CLf.UP.,g_e>/4F(YdE>4C/;;0@a@dbJ@E;4XM9NY63H
V^7RBU(7[S+9A)A^2(LTF8QcG=@NUf,AWLF+SX1Z[2.I8;E70eS1/,JfJ1KDC(K.
.>T3J;V-?FDgG>@2;NP]UUQZ3E/B-QHbS&N[^0S)53CaMTJ=>WD1^\9SS?R1I1;e
RAV5:@e?bAHNWZ7A4ILUG6fWX)/YZ2MYKRB1c2,:@XedUIF3;6O<KcOdGV@T0^;=
3KP8JLY:6YfaR(N\^ac6IL_Zgc[FA(e:b@2Y,>2=.ZDP^S)XXT)):PgLHH217&F3
BVU/EY/\f->&R3Ab6W61D075B&^(+=5>)b:cc:2G\1>aT[Gg2VIgPV6^d8VfVNQ(
Y:6.,OMV=ZODHV&]SNCU/^Ec(1^KcfEJa;OC#.7B:f&;.K7&>I,edB5=HeUNH+/_
S2(F[1+?]#J_MACd/U,@\@;16Y;d+XD5#I]T)A1g.RedC&YfZ+Z79AK[=C6TA8#7
V\_F?@f\&^H[,dcR#:DeLca_GWdf<@&>DV\>?SO2LFP+(<?cJ;g;4#a?KBd_;dCX
;S\N8I7UR5IcA=I3YdT-2/IDd1_e/C:/WF/8,3g4P&7=K\L5POe3=80CTbJ^Z)+W
@R\>Zf3M\7de@LVKcg<-KV;-K:J/BD]3&G#.2J8aXeZPY?90_M(KTA#)7+VO89<f
<NMJ;W2L[aQ:I:XbS^WY_K^,-XL0^Z)d,Q([ILIJ5L3UBIVW3@UcTKa4#R,]Y/\^
8HWb61T/eAWd)V.<9K@M4?ODWd+cTO]\=3bZ@9TA2BI[Y?#.ZNJ3bSffD\/C&KS#
1Z/9dIGLJgdJQI)bLHHG-Z88/^f2(^?JMM_dRV</.XN6VM5D(1M3@]RE=cI]77e@
Qd=IQO>b/+@L3N&YfU2Q34H)]@YBSG0QOLN[,N5[eLTZE.W?CcfE6(5YdXa#GQL^
:E(+LR82Z^452[R_FK48VF?D&S29/FfR<cL70_>8@be):X4FZe_2HPCL(]Y:;5=?
Ue7UOV?@U02S]AUa;BTdACW(a(g881GJf\6QF/=LFg3DSJ9LB,W1-8#>f-aM]6/U
2O2g);.@JcOVUa8AGXNKVI:IO95X:.a\PL^Jg(Z\]cK;XTM98a?=1J6MP]0&2OE?
M,\/:I:C=JDOdT3ZBGIJY[^\/OD:-FC6&#J)@U(^c?A-5X5JD-WQ:^/G2g<JdZ-4
,Z7T)GCfMZI/7J1P_3L\W++M]a]+NZ=<Y=DB:;>U6aK9d],OFded<K)V3R(5PUNR
1O1d,3P@0<#E/=XYD3VA>M7&J5BSREQAH_HYc(Od_7>Z@:FC\>)9.3_92Jf.V][1
-T]9.c4;2#DQKIJ&5JU-WJ#RI<H.(A@_Dc7_-AY7YCSd@D-1gO<#1gSe;F))P)S#
.)SGI\HY:JPd0BVFd/WM/GI/L9U-TfJ>eVf090c81+1^-:e?PS#D#@QCR#LCa&Y_
CG7.RSB]R>AIF?FTd(8:2;f4&4d6f5Sg04J)Ab9<91N,c^E19Gfca]:a/X>8BHgA
8V0?VJeYDd<B5-&4RK?eS3d+.ZK9E>ebXOJI+cR1K7T?&Z2/bgW[9/I\P#\@>e&T
^VO1B0RW45TGL-DC<&Q(^:UDSB:P=F.->/F2\]\>VR?XKOB8)#2+=\D3/B)44fg?
f):XQHPVff-XEU)f\EA77&O6(IH4,672Dc6O/UOW\f<1^Y,D70dE6,L#[1UJN8^9
E)5gg?eQ3#E8gc+IW;f\3[c-=TIZL^;QBe0Lf:?baVMJ_:6:]X^Z_>d(&Z4F2U#5
ae-32Pc;L9+8P<=1YRUP>X_QDGFGZ9#fP0I>A[604</9/Gde@4HbbSdFa&IVD=Jc
)ZZ]3c-=D@[R2=YT_MggS-E20ca(@V:2G1YUL;Ed.Z@Q,&ZO1V:.26X@NfO:Ve,T
7&>fVC;,@5=cJ]6TRY.D9/;?MK7D#RSJbN2ZM3U1:41Q2],;LAc>(B1CffW/Q4c;
IP119_a<K?U6UPgc<-5afNT\B?342bUP1X():<,C(=@5G=&Sf^0aTY8^F.gC1&,5
f36^.1K[/P@+R^dgbC@Zf5(E/f<c>DF(g[)]@^OQ-ZSBW=;+V8U&[Y4+3KYH\<]g
NIU,1E;Qd9Z4-956V)N7:@^,ON)RdYYB=e8^SZ6J<\U2\?f>L2E;T20Z/^LeB/-&
I4S_?5^^1W:QSfb,IdQV:WZ(f.?AN-:CP6IHMLX(L<g3B=XC<M(>4d5fR2?Hf^]@
)I>\d/+:SW\aES6@Y#_4WT0?L#0REfdWcD93Rd^PD+Z[8.g)cHAYM3N8X#[[Z/;#
/?V=SX_C7<bdA[(/)-.99L0RgSB?KYVR4CZ?H=95eQ_1DJ,6U.XQJ)R^(?Fd6LJ[
ZZ?)AdL7.MUEDJH\.+Z;3JA5LA\b=L0BX(a8_8.B];O>OJ^6=RbM\0+IbM-cT2ab
I.;UHDRO12#-H0MH5N).HPIOg#?RNH&fW@2\[7\g4af\N68dF&aPOJ3;K99CfV7_
2.4eJ1]OF]HIT.I&FH\&2E\KL\GF/G4VSd#U&;1[&b-3^>9DS:(9Q,=7dF^Y&ad-
#\4=IC;Vdge4#-]BETOI2>QLI8J1U57c0G7K4fEHeF>;I_XD-G<+/68;&O4]^BS@
AC&e]UWMadgF36.Qg15<==M;L6,<aCNZ=DS\f1f7]Y^:)fa@TFTCMMIgJSaFcPAU
XTGg,=W9ITA1DKC>)46_#VdSID_UFcgJTb]FN=CB]b.U]X[N6V@&JJW8YI.0fb)N
&MEKV/FXQAP]&Cc/I;&G=6#??M[Ee+MUYF2-S@]1F[X/;SVe-[:Z8EA+F2:YFE4N
T^dQZdQRI7_Mf,3VIBP,_1M>.;)7KPIKZ0_@?\[_gN,?]^6T4+QVTHL(aJ;b0;e6
+-Q#eJ93+f]Z:#E.RYIAf-.H18>X7XBEX6GB)CYLNga(Lc4+YgK=M00=,DJ;&aA&
6ES0Fc>E3bE-YObg<L)bR@>A2C,;09J_.W:Q(_YcSeA&e:Q[WC8-?g,c-N<RUVC5
7bL7#aWPaAX87^aXYQ3NH+U5UKTa1-BMP>cKJPOF5><;HVN.3f(UM#H+?2>9:_E?
5K#\?+=c;8-E1M)fLg[,3dHe.\4AFKO:F9Q>6gP\dR2QDZ+J0;J=RPSZ=19<O03\
A7a8e/COd2?Ia&7fc#K[KOZ,(+7Y8F/<9.0SYZaJ^fb,YGI0LV@6:)_7U_-MCL1#
,fFe\CPe3dKLa/FXQG(IO@,&V\:R&8V+^T=^K8EX3gf<N<<bSLM5Uc?B)[^d_L4(
5acb7BU0<Q7CQB.cA5)C(T,[].3A[:6-aG82(e95<9Wb5(P((K/C=O+UIg+>_KGK
W^;+^F3A8:#XV)[;:N+8O[<7UAB(6bIQaHP1LeNLP60W+J,4.P]#e3XMK,.;I=g5
6N&Rd+U>1T0@bY;ROE_44>a#Ja+cGV4@(.^\,D3_GEH<-MPZVdc3E#.Z_K4F<H??
Y^K>0=S2;H9/<P1ADfKMGf1T@9dPK0,CD#;6]N#=K?=?Q<W0OdcE[33+ff84g59#
:X^d7dF1H,C+)7U59UL]3aHJ4W/,+gC;]2<H;ZK8XXe^2c3&C29<_F3FM,?LLFGC
0_=H=<_8V]&U#bR5a5):WE>)BIP<a\J<:YQaF-]JPFIBdVBBOP.7>.1eUDR8JYN>
/ZUB7XM6,?>.<cU6/Bg3b9f](G0TV&_FRWH)7-HY[^&,cRf>/4cJ4,OS8eD4eO4]
CPFE4eYH.fLX7H2,\Aa4ZXF4KBZC&f3?I]1SZ8JPH5)gJE)UH,g<ICZ;2NbERbF#
NWXK[DE?[a26MgDRLYX9A;<f[E8RO1RbC\-GY^)/:WAA4DfJDB7V57S7W#-/0,G/
2RX]L[&JY9,WI\KF6=SV&8E>6HAf#g9;BD7;&_.b6(g90WDgSLA\F0)DT8?JU@aK
@S=WKF)YI&[AOg&LML>H[&HCE(CD(-0fK27?)IYU9?&a;8N<d@H(eR]Fg61/e6@M
H(1WG);a5_)O2XJaD_5A^-fW]d2YPf]S<:CP?MZ/4JKSGUY(PBbG9gK8KaN0&#_S
\HLFVO>/]U5;9<@,M9[0,_[WODU5/G>gJ;SNO6A\UX[0;b(EJbM@4E6/JP6Y.ZbZ
J<<7H9b((aKEZ@Qa?O9([+c[Z/AYH@V>dT4F&J:(6GQ;4a[B\4gf/2Y?\+IP5gQV
<dAdQbZ@EF5a:U5&286>/Q?>Ce_7a0GO1EB=FNF9-Ha>K3eL_+#&EIN7bZ]4a)66
1PIU>V2N;&a]]f-M(W49D#OXUX8:NV8)A(.bDYA^a4C._M2MLg(eZ&(>Xde[/??a
cJM/)RYL+<8BM&#\FI\\+=+;D74WC48cTFdQECC]B>8^O7ILTB&U/&+K[9HNB0=O
E/e,T)714/=\6-QD\-:M(-GRVY\b5gX4JR45Nd=S]\IZZ?ce5fH=YCeP;]0aBPB)
eZ;LZW,Vb#gTB22C-S<7]<5UNK-d+,Y3#1SQ.N6c,g+\B/.):8EA^SGf\f:?:A=8
2C[YK(X/::f.]T^YgF2L&WeM&Q0+IW+P@W>[E9RQ]Z_I<6,46W\KdAcQ__S5^F5J
:R70b^\,?9,H);<Z16BP-MeII@L_F\6V?NMa&^MYUXRaF[[NRIJB-6LCeBNQc&dM
fb<@&ZRg=cb>+LgN?#,#=D5K/EVTTc,7f+_94Q;U-+@<N6LL7eBY^PaG9+;\11P)
Pd+M[_/HgFIe6NL1/F^bR@57/7:HW8FU=T2L:H]1T-FVWB(F+V(.<<;[]J.#2G+Q
7aN,7\SgGaK?a>ef1?[7e+[P4T<ea5:AFR;4N3I0^I8AD<-M3f(46>3X86_,3AMa
5&DcYG.L@K[X1];]/3WOg(DC<eNKX.a[UKMR4+6(:RXXc0Z-V.JaU4H.HF;:AO)2
P&.E\g\\2-b6R.2d[3L\L8WB+/b&WX,;?7f_E+N>ECUJZSG[7[]FaIJ9b.A97d,>
&_G0>U](PbMP@5WBLAAJ0^f6Xe^eDd-I;IC>A>E/##05a(F/=?8X]1-:O\X[edCN
UBT+G_1;JI]]Kg:.#baWF(>c)-4\C2/N^2V<0cO:b-.[ZK50I8QA?\c,/NT]->DD
=\#6<RVEG5->C>Ab\W@06N9)M1GD^MX;#AUHSH:I</DH9CR/]aFJfeH_b6IOL1c0
BLGE(4>BE@a8-\W<(>]=VG95?3?2,8aF.=^>]Q5_F\P4LDKK\7e+WaM3&=&U6+?,
SgJN#WFUMIL<V>cNK-OV0GANa_G=<0;&g0OG?+IIV0E:T7;?4?TbHIT@1X@PR_f^
4.aPKOQ<9UMAOg]0[)]fCSYT?eEROFLbND1g?&FGHI9_T7-7Q&EWab[16+#>0f5<
GN.5,T8?8&Y@C3aKS:MdRB]8Y^acWQfTYM9\a0G3R=Jf:DFa1dC^FN\PCd((;SG&
YSN4OINTNB=.40JMg1PBPa1cRVGY4#=Eb1E>6A.A\V;N\7MQKJa:Q1D0V.fJ&QT?
^]DXTFJ>eXL=Dg/5;)DKXdJWK(a?[#5ESP?(U[BP89RB[&bTE3B\,f(]@.=N2^)I
0M&7Ub1F4D[J?M&8d@6)BADH>H)AH>E3:@H?UMeJLN6M_Q+9P_=C9@_UEBe5FFT#
.cT^86G]\2=S/BBU\U)GLbc(eKfNEf:MKGXXe_f]bGIE^I0g.Z63AGG1I7K:,?ab
N4#I1U<W<SbAP[G0b7ET58TCNU/9aC;V&Y4Ne6JHOIAQdH8/KaWSJ,#0?MTO,<?7
7[7M+/9]c]f[Db5.AO6)KZ@3-3Z1Xb^DJ(I+/9g+&^=A.U5)ee-b@Jg2K;d[#-2b
gNR+-@@C]I1D/]VB4JP)b),13PSJ2\(+KQVe&cX5I@d(3TPS^\>>S,YYb_Xba4a?
@9\e/HLXEVSM(N=\Wg1J(:cfY.cW,]U[>)b7KD?Hb(e_Q;HHF01M@aX,aAc]RHFT
:6:B8GP9RcY+^Z+:b(VN:7CE1ZAVE5g=GUae6O&DED#99#VD=4^4Yg1e\88>V2PB
TPP5dYg-?M[8FPEeP>.YN1A(D?_0COF0;MCQ]H^UIf1F?,^CIBG_Z4/SH=b7cb(F
B7[SBd,R:M+Z7\AWIQ,X=-O,.&\D.>:Y232GB8@P:>ARb./+8T[P/,Ze80WL(NR^
S;<c,XA+8-](SBBY^ZL\1_^M.KGLPg,_3PY^9>6X+,9;:OV_F_<g>I51RH,RQ4c]
aW#>fPPW()2G8Icc7:.,VeUA,#PCg<f#-.X_YW^:\TaORd&A;:M_:/UFL=+^HFNE
(0>/\Uag8?N2)UP:4?@S3?a^:3P\/U-_,:+-YeJCZTQIgELR?S,9)_B3J:<:\4-b
KT)##f<4W/5Z:dgcOXVOeJZA2_#E1W5U<:^R]JG#WF;EU??B@Q4.ZVS76F9[1FU?
N-GB)>H9_age+77eL3ECc<agT3VE,4^@4^OLE&=C,4]RGV+eF26+L]93Ag]d;(&#
gN[.5P??T=Cde7OH;(/A_TUY;]LgRVEbb@+9GYAb=cBHL0Ff_OVR[RP](Y4OW5]X
5)AKMTF_,B44,:Yd:fG;]RQ4N\c(AbT/<Tffga&8JbAJ^C[G6T05>0Na5<Y0bEUF
CCK(Q+F:D:,gBC&>H#2P:.+[=83@^ScH7T5c);AH]VVg[Y8M+M\?^EMYW:MA6f<;
FD&90E6PeCSO^D@H,\D.K@,Q+Z8eQ0.N,-THQ<)NG8C2;:OKYE7TS2D-^?Q[a6C7
O5G;fZ)-=?)NPD_fWJ=2H=\X(]&ES>1/Qc>FdE4e2G:^5??9;JO]+]Z>E,(^e_P.
.^DP+CCFQBeUN9&JNaT&G7PH0;+D3=gddLI:aO2PT<APB&Tb11J6f6SB416=K&1_
5fP4&<<#[:@?&K_ZGXS#Wc\-ZW93e(=.?(?CF_X\bdBA)D?UX+1aQ?/8G@_L0g/A
>Ha3XV,\)K89W]I&HM47T#Xa-f7GK@1aHKB;VC?U:>@G_32gE4_\T0D3RNZ45O+b
K2f,VBTA?4b_dQEPC2.DU^P;T9e#V,R6\+U^eJIHKDX^8RGIL3>8HYdVV#a9;DXT
P/-(JF7-)-QZETVSfbf=-O)8;._U,ER:B_._8I>Ud2H8PE@@CS3TcdJPW#4,3QaM
JEJBPNd)T::eeV&FCSaR&bbU-+31;L.)FXC;TU:?:1>T0PN\bV;KAf8DJL6D?V^=
VBGgM(ONRO&.RWaF;N6D_Q:K[CF@#,NY(>FX9VSVDfJ0bIXCQ#S6R1S6FBe,DL?_
TYT[JK59Jg1<;)V,LNLbOOAFRf7KX,GM=QWQ]R+O<6DaGRT34aL0D?(E=&=R7FRI
VQ&,3g^M[H;T1f+<#[W/b47\#acD7<;a:/2H@)0aaR9KTB5K2,O^YK+I.7SX2=(O
N9M0IS)=7U<Q)][PD)332>:9\]agF_c=0aK4b53)Y89B4@)K#)]>5.G.6N>;fd\G
LU09T5ZPG(06a;:SX=V]-S0RBKOVZ+1UX&Q8(9AJS46]=FNXI8^NN=#8:?WcXe&3
M24c2QGa0,V-S.6-I&K8bGSgVXfVBLA7B>E38T]6URf3</;5L_F([1(_cOU\F/4<
1NL8Q[fPfX#K6ga(DDI,0,Ac--X]^OgS<YOeJ;2\F(f9T<B]]a4J#HOAO+VS+H=^
_)EF9MBJbK4NIT_GMe_9@7].FEI0D)[_:^Za)HN=]&]U:+g0]WQRC_dPQf7Cc3W<
RSF4>\>=01Xb+0T?=O;4_cQ)4+\RQg[>cc=M4WVaHOZaWCIWe:U/3aOWLe99^c9Z
UFeWe\I3gUJ-DYf_RL]f:cS6\RHZ:G#PaRBW/aR5PbWQaZbbb.@;,/-?2c7;[,dO
UK&PU8^eS(@,?dX:bRC7+Hb1GNIaHLA5_PDdY6N=+cG0E\H,=F:05,#:2b,=3Y0M
9QOT>#2=T5)3_5?b<H?a7)\Z1Ea_CUZA0L@FJU2V1.90:YEe4FT?WV@2]7,;:<J7
@Ue?_BEXN-9BTf(d@1g2K,OU#f-R2.fDFNZSH)87>c:E>Yf\7#,IZ9\)UD]]&S@B
d1+\?(FW?FA5)dQL:,5eZI6E6PVWH+&.F+KGFJU.<2c84c2[ZZKg^JAgD:7gVK^7
Xfd#9OLg^57HA.cG_=,<-NFYeC^)EeCba[/W)?+(,8[66dZb0Q?5c+5Z6EX)aSgI
&Z/FB87^RG:_E9VdWFH/eI57NTE)=/#HSIUA&I9+ICU)X#PW,VB(CFX#B+GRAbbV
_GO^dNO;NPTT\9QNS;_C)B[gM>RL:>A)5bb8cNLd>96RF4C2NSJG72dBZB@@REba
a#ZLS0a9R3Y=(U+-<0.ad)XJFBV\TcHdR^H^CVMZa?34(^9K,2GSSM6HBgWJ_?[6
#bI;OD<I>Fcd@N,+efHHZ?IV1QESb.7UYf)(>LHCF-4-0XC./T;MVS4Z<IfXX)ZB
6UB&_+bOd_#I#S22<9TQV?7B6?R2_VXF>DZ>L4@dgeY=OIR]?&<f-.#gd-b9BO1:
3g9.?f2W?&=I2Z@)dW47@K;A<7[,:_fV<NKGN,bFR&d0U;VWF=+Z(4M/8,SM=6^5
L]:R4,a\CTKbS?G9#:LRd:V5NVYC=WHcIa=LI.H^:]:+-^R[[0ZY=:a/0E//P7..
b-\7R#D5?eSZ7((1>.cb-3DIQ]eVE6Lc\I/a_7LeH6AHe->;5V)OX.3Zc=/0F7F:
-^^+K<MKKHSW#S9/_@c8Y+;0KLf-^RG+)0,X#MKN(0&2#DU_0[<J50+fX\_97W<5
1FNDPe@)>:48OJd_UfYDQGBW:F^H]QN-5_GEEW)/87@<OFX4T=N2X9GUD.0[M<MV
X+-HLZY@SRcP?-D#]_QIUOg1][3=_5a1\3-MIDQLe@^8-+XIRGRB-X]d[8EcM@FB
Q.)f5\5LdYcN9JAA>AL9F4?dC?[(K)Y+MOd.+EILG<3WUf_X8H9ZKGcDKb9[V;b0
TTF0Ag)\gX#+=#ed6(^3]_,JFDKd\378FIID93M=N9=?Mge<47V9YXgU0TM(&D2\
)&IV_LL&&(^JH>-FFG^WXg:F>GFNV;aKf?JfQ9PI]NB,+WMAaEbe;;G314/944IV
I986(8WK4K=D7Se=;U5#,TOQZOT=MLDcIS6)?ABaA/I940;93CdO[>1AZ^N_f1Re
;:/K(H/23Cd,<AS=8:GQ0_D/dbJ-dcS_e>B)Y_M1d@K>7@QM@dGf592fNVT,eZ6<
_<da9^TDU;Y+_?+OdEJIG+HEJDPH;^da_fCUM_KXW:8-gcC,-#:-(H3[^;cg#<#U
U2LM/V1V\gXL[N-TI\[X>#,SX+Y<Sc?E+/(DAP+0g&.EMG8M-MO[DHXF3-[?2R)O
LWUGD3KAJDYaA<gDRCG73-JZABMY;V7^CK[La)c(:O,-fV+]D@06\++SL?44C49.
WN?<LYBPW2VE^JE#KN?dd3eGUJV>6)\L=6.)UA+_6OLGYZC^PZCYXY>]J<F?,:AR
ed+b12?24B-;&:0bUTBWW@XP8F=<?BYMCNdfgY[ddU&O@3;3]H#PJA@57/c9)b<C
^G+66I#YXF:\CB/#NDF_DQKfDY0N_@#:f>>7J,ZP#V>SDJ\YMB9?Le@1QVEe&3U:
\K]Sc^^;1<=@Vc@6F#JV[a#+VHI].1N;9T<dC;R-MP4&.P@MHObFaGFc&G/M]b?-
#FJK/927]&eB<OH5KII)VW)#;CXRA0#,IO#D=(1I@P;6c?)YM,c=0DB_#GK>0b9Y
dGEW<Ye9S?P]X1NO:33Ibf?2b8GE0P6G@]8::Bd,<9/9TSZ+0G5BKEVNaSf&K38,
VCVb.AaQ1&GG\VL67A6cU\/MeNa5]P@E_OJG7g(OHS:W.K43EUFS\(H+AfSB2SVe
ceKISZ[>X\N7ca2e&&NXM2c1M1XK1B()+:(2INZaCaH^BR8BEafg-6@eR7#M]6J.
9&<AI9ZEE=8c5XA=Y5eY]RIMa?Sd_/M2O(E/de9_)3Ta;DM=Cf24=FeQK&O3_.XH
8I7FM;WH7]E&fd[4W-N?@7Mb1+IOggQUe(-K5OgWP+1LOX@3A2?(P>62O#OQT_,&
3>,/5?JD#c+RH0VN,f,OS-_VeJ]WY)bd;&aY=YO&=E8ID8,LW2G/gO6)7b8O\7;2
M/45B?7d.ZF-<[J.HQ68V5.VVM/(YdTY/KNg?cJ7Z+L[eX#>N4=&Ob;G(8XW8<M_
T2.X57Z<1GUQ7.+3HA5:B]b+F=e:f17dPA6Q/.Jg[FUf/,+>Q&Z3;6XI5bc0[LGf
RC6;gL=&^eT[JYF2g4?7H-MUI?ALfLK:0=EQD?:J1K1)P#SJW^[X:YRQ^c3(5-4@
gN0[\/\.J9c06(daWA(?628EAad@:,]^NXd9b<NK=CVN2R5+B^:Yc3_QT<Te\2=.
#VZf@c>E5Ke-N2@_<_gC)eY^AM-JBe[=[C9+1SLD^OX&8eRBN4]U3;)JN=8R_UZJ
;6K]]^Y<\7M#+TC1W2EFR#b,E4f?;XC<SE]AX<M9QD:aA1\cNX@8-AW>I;-[HP-@
1P>0\1IM+>DC.&H];FY[BWeZeLFGbQ11IHMc23_g>H42cb5Hdd]+^aXFQ=:3Va,H
,MN)HQF##D)2:WS?X,Y\)CH?4GJU[OKAM5K\HAP_<FO<LeVR;L=<HQgKUH&,Z\>c
<(Q:2YQCO@WK./d5^\]IX[:O>1/\(c,c4,1R(5\8MR:Y#I3(M(>QU4]?DVZNB_e3
OaB1a6UY<+e[.NC]JW.VcR3BF+ZSYeNcVbAc0B;K?IS.(S1KM1=8U;8V>7Hc)L+]
E3Y?^M+]53UF(1Rba02=UHgV(1EDcQH_;_9bJC.X@W7RITCf[(B[73Oba)SZ.\^L
MO/HH]b)BbV3>Z@bM3+]ZX0/G>QB4ZgNg]/)C-Ve[\D83A2C:H?3=OI_7H&0TW^M
VX0/7[b,Q=cgRb6?&QB:(K:6\)3U55W:a]KI5:HPZ^Xb,ZHASccVJQ=N?Qe7HOdC
Ia)83b:2PMfJJP3<P-=)&^6--;>T(K4T,_JCERJK#0=9]N6C[9+BfE+)LURM6Z9@
&__X^JC9&J<]SQI)9Rc<5f1=26(3IK2,(H6V(K+()SI\+fK5X(G5LORJM<(PL0V]
;gQ(XK>dTLO_FPRQae]QgXgd=GRZSXRO(=;71;>0Za:E]BNbK+=E]ab@d6d[.VdU
NR];P[32a8PfL3R:@A@JHL<HMKS&_dJ<VHMf),c7.7ZYNX3cd\-VY3B?F)48&:E3
cH<Wa_<K-)OX;Q96EbAGNDVASRdI)BH>K_8B1R_<eO^#WLTAWKDfSJ1a]K1BUXVb
CDXS6LLIbQU,9^@FS2e97X@37:^&dbL.6^FVJ^H7&Z.,VGI41G/FH:B,@Mg\AT/X
MH=A,PW.+<1(^B7:]XC658-.eK_I2SFM3;R&LXWa-g+EG_<.5<G/=(a2E(0IWLR.
S/TL3(VAa5H3XRY+F[K3#[A6(O8_^e?F-3-70>,/@UYB^KaEK,PI.a]TI;JZf3)>
MM,7_V0^&6LQZ8Q7a3O<]T&a?8a=:8,McQXYU7HG(3ELF#6E/V\2T]aG1?^64(:,
W96V#/QI5?aDee@DT6D7_WA<Ae[,P+]K2B2)1+G#2(.HABL&O2HSC-IB;R]PMRaC
2]B7M)7=#BD8LPY3AS,#Pa9\#TT9CGdUdB+?e237]F-]-^]>Y:BdYAU\7DEadY=I
JN<+[<@/Z&b2XR&;I_YMaEN,(>4gWIDSX7BE/=TH?UD<cTgKY_<&WAN)[ST-8_d^
RI)]#5P1dCZGO(1FD.HLIS)RR?P&C\5X5<=@X89^M1BORO_W0GTNXEM#edN1#a\3
&/dL/B/\-:WK_a^ML69g#\2EPd[XbH)5g[HaUJ<805+I.;)1;#IH5B;_/McKS4>]
?GA<E>g3JOR1FfJO()^d6(>Ag7^Q)J6TP09YLJDS6BQU]_>/gUS2H+J7(e#7F8A@
+,R_I4bK8a7U?.168NNUX1+)(b(fd:)[TV2Y+XAQ).+Tae23:(W;QC)^CDQ1Md_?
3d[UFe<&T=>7S;2MXUOeT23Nb-=E:Z,dC-&0X09c;_)K9D\<PcZfML5>:I_J6-N[
L7EaNVP1W0b5UgG4ICeeDG)>,8=4J,B/#We:Pc+\>bQTH-&,PMQBCbOOLaZ4abUd
dZ>ZI6)1V=,Uf+=J4G@Y-55_+H)cf8OM[Jg_)A-B]LAN0L#1)5JB4U[HQ#9IgI3H
#Y=fFEX-CWFV^U2Q#X=S7@&7::(P@J78RL/UcaCObLU3JL:10gL6#9^X^P(O/MaJ
:D>+Q;(2gY.c^]4+/@0HQ@Fe#L:d0EQRVZ)I+1OD:3+J-U:Ra4^fNE_a-KZbgccG
1A_6gd3W)S)g](.KQf_6J032Bc30P39T(;\:H4cR.BbMDedAU]>8bLB##8,]\[eI
NN9GDcCR4#M5@K#3d=aNY2/)IX2Ce^CC2^\@6<]F1aVAa<I6\(K@U6febV6?@D\6
E^aZEQ7[RE;<K<G+;Y>AFWb#UN02CG=BT#L\)BK#f&=:13TL:]5BdK.CW,58a?+G
d-8,:Af.F<;M]#?Wc&=8BY3&PPZ00VN1WO=a^>?<W=6,UYa1g0dW[8e)N41C?NXD
_6&V^TL]#[P3Rc#:LIHJ?NOad]gcA+ZWE?8.Z3Q?+K&ZfMX)HP(f+f2;\GQ)[)N:
LN^_L@:AI#24KeY_&<23Qg3152g+AYcYYgS9Z48R\bXS-@2]0:URJL2=A9EVa(9b
fVPUJ:MO]Lg1O,&L7gBT)1JM(Z:c@=:Nbag-VgPdO(-WWID_Iefb<P4R2\JF8NP[
&EV7-&Tg[,R+_@dI-U^JUMW=&b]D+)+;K4C0H_MG:K/eQDB>Sa@,V@+]BGF^O6a3
f3=K>?L.FL@32MQ99@5_SX68/C]K.;W.<dJH_T;8[.M&LI91T?Y.+?FG&<M3XD.Z
Vd+VcVJdE?:X-BZPN-ZRE4b:]gBE3=>#H;<0+Ma1J;R34KCK3+8(c;9PVbfWFB1V
c1JOd-JYJ/JY+UBK>::&f.D-LX+>_^G-,,,E&XBI=/?8?2Hg10RK2;c1BC3eg5#(
BP]fL3@GGbP1J1_-e2#=U^ECX]8[OgcW_53@)\2LPcNDeR;g8JHfJN#R654\.99J
P<A]=OV4^2-NA2<Y-1J+H6OMK@/+@US\R_@7B6UFK16.1W+4Q)Q=gP4V7\1WUW?Y
SYH8Rd^a()cEd.PT.AN=Q@Y.72QUI>T_(^e0@U?Z;(KZ/OdX6e8c#>BN^&=W2W=3
JPHDO4;7IeJAc6JB0Gf-dd&D:fT,6T[3,Aa#[]EY9A?,aZ,[:;E\[5N.@9XL4C(B
KK==MB[VMc[\d?FWEOD,X&(WC4A6a6_LSF&L\CDCV1BQQU?/GYG23YQM+7\Jd1\A
U/7VB;W)1-:4V?GLLPUVY;6VA>CZgY&a_):g@0c^E<STL2CCGd]V5g)B(447c;-B
=-WE.A5Qe/[gJf2gMgDXM;WYE]Q:[eRG2KHW#=f25:4cfA7NZNH7FX\WZ1Z80aO7
,<2]N/ZSXYbGY;BDJ>VY^d8\beZRf=H4],>7KZ-d(8A(?E^APJ0(]W3^[_;9>A[e
S8RFJf?^1P)D1@+^)V<XWBV/^b<&Qf[]D8_aUJ(3)Ka+L(2P^bNKM^?d:;^C[KS@
E(,IagJB/VWTUK;6DH6,&Sd+I@>HT@N7YZQW&C51(88N6JdeXA2_D#ScH+L?Q\(b
>/N#+.W8A/LKV#[-JDCJO.[5cG3RNdceI4_J(fD.O5A[TL\0UCQTa38AU#,D&M(:
;d\(1#CdH(#Y?CI-JWDeRI[/C4aa8K+;dQR0-AJF^46G,[XLL^Da94_R.,W1_6,<
-ZTU42CJ?5/C/8ID508B-Tf5C9W4-7=a;,K:34(H<-V/,S]?O,gX)CX/;Of-a>8d
[RXI)^cI;SU&DGZV8.L;XaK>H6ATdS168PQ(3#/7O(Vf<OJTd=@6U_/WX?LFW3UQ
ID8E.RWYDLCYDQ..dgN<SWce2D>cJff[+\d>HI42RV3BEC.[;/b-g#6V5[gGSgH:
.5.K#<Gf?#Zf,c2DXd+0T:N@GA@J:/fZ^fM@NYCH[W?1HK//S2G\.UI/0U6eGXWW
L_/GV(/K?@+8[FMS<HF6J\2G]6Ca1HGca.X(8X#b<\V[JYC=RZMM9:NY[55T#ZG5
/TJfY5RKE.a6Y94E58TZ?Zf.W/IH[C8=O)6(BFH+HIC>ea9S?.4@)1_6LRXJ<?M0
5IRT#T.T#&QeVEHB&@HM\F9bGZ@5FBF/8SP/&fO:AdZKK\+XOE7@C8,R:=+=V1/N
FCTOI?dOf[817NNDRX)[@,)#^/Wf[BZ@@9XQg5R@?)W)@_V7[MI4e^]5EZ-9:V&P
M^=8X=U@1>;.WH0/A9;/6/-2=0dZd8&YTW8-P2-SfO9KMMVHC^J_D4&0TBVVX<-&
6?S.,Z7YC9bcG\g-DGcU[<C;(<\aOb2>9E=Y8cJZYCMAS&OQ7G2T63IA1NJVT(_@
;d1.AQ8K_7B]0[bS(3-g[UK75GXdbROfdZ1f1\5UI36eWX=)>UG,=6ILgdY2UL9>
DaTTa0-1YIdK(1Tf1),@dI@9;LP-gHC#>eLNASI8[2^a&f2-SSJ;R0#=ISG>=?3>
.32(D:_fa9J:)/ZQD,<@RT+.K70=,4GXK7R^4>\F3c4VgG,We@9J<7EB;f^(YUMb
TMJ&TN5K?Y;O=I868RY@7XR?YATLJ^:\)-6<?[CGWY_4R(([)1g>D8?a?AG/0XV0
9=UbVY,KNEUDCY:-CO<VCYQeFDDg=TM(MTU9We1RUafd;V\IE\K]>U294\KZcVS,
MaSZX21&,dg57@ZTM:DVb_YX_Y?Cff?PQ>SXT18ag6_Zb&W)B[5=0K@1?AeB.J5&
KF/GB#7/]2]G<EF689\]T_EgXYA/T5aYe0<?CKE^6;3f^7468ReO_<\^_P#O?c1-
_JPE7cZZ7eFF7K\K0<6G9H^8?49)]V17>F=<0B_Q3N-T(YWgT:d[2^>A6BIe)^PC
SE.ZGDUBQ06IXA]#GME_=I@fDOT;\2&/QD&GaQX]fOX6E;0GcV]Z1;#DYK?b@,cF
SC]NO9T8:Y+6[AC8\PgE-L.8#c9/;)b:QR.[,D+eNO<O(D,8\ZC:#6YB]C^g4gVT
b&3D_OU/O-_<Y/2bR4MN:GdL+c+Q;PVP^V=0,3_Z)^b\eBV7aSF]b>.b#8.E3gf=
U076GE+<@)G&@Bde6KdB^:XE9WAI1VeZ2a)3XU;Z^UTZ_+<JcegP,KDCU/?V^ba0
.?NE_268TIMSL09-f.+[1:P37\JKZ<gZ]GN)\a7-H9=LbJSI73f<d(C6g/,)NC>c
Z&d1W?H\KMgegOU,YNR86,JO>Z#,<Z9c,;-7=b,UTGR\gVNCO5+5A=<&O=9NF2V^
QET7g\QNA63&&#QVPJGTQdEA#A895YLF3=9PB;XSeX)a][bK:b.G_EF8&eCZ88GO
I3Pa]NR&N\N(MA&\8X(^b+S(+0LR<^\MCRY5#=eK;_/#SVU_2?2YAF2-N994,ED0
X#\?J-1LK2ZNdJbP;J70=S(\>M)#+_Y]@]HP252fF9:)Ia#NI;96>c7R\a02eO1>
]P5)0(/(VQTN_NGBa(HRKg/Ag7D7,FAdf:>-BGXg=>[fZ2TT413dfHaE^e;)c,5H
7N6#7^#2IbJd>@2\Y7<.X&g/9EdIW+5)&-4H#5XZ=EeREF6O:1a=1:AM.MF97=>_
@_T(9#HW+,aXXKLdOB@R]V&1?)ABG5=;M?3Ua(SM_a1-4JcZ92L^HOP<1,.GdFUX
9.&P\]2Cb4dW1T(5LCH]>V##Y?;V8FZG.]PVPA@2L6HaI9fPFN9?XE0RC(23-@e2
T9Ie[C=KdJTK0+gOG>L@LHS=I1D:WJ=Q#7UU8&(2g0FJ^8KR@_7L8M47C66NNS4>
EKO\gS?1QN2Y)b3JcLR<<83]SH3F)WMO6^,WO,bK+0IWHf0,XZg_=9H9K_9_SMXA
YEI:LMO\BGL..gR,feaXe5OE2+CQ.C5B.^KI0f_eC@Wd2,cL.?5W<X)QaAf9I.\J
=K&\0OeS3&IAR(D7&7baLCc.YDN/=#dbDC^LI<MgIb+gB4Ga-TN^S3UMSM<_bA-b
K.dIBWH>5S5D6FZ8E>:-HaN^b6J-:Q+_+,_@Q,N,fX<E>9KI.Ab^Z5@DZ94UNZaY
9.-Y@cE/QYE_2D)E4FB3#[[SUEc@=WXL;H[KU^8NVQ,/Lda30B4\N+Cd##:G7W?1
3/A5&deg>=&..NXEQ)7+K=R<YTT2bb,AA/F78FF5>CN7K:/8IK7-,)]/1b9008#=
8g@RPC3eYI3R_378[1_14BcB8X_M\G#5CUBC>^;dZU\K7.=V>e1#U+SX.XT.R1(]
g=^_4EeX207DF49-\F/>:K9R(cV9.:JJgA9&MaaI:>;#NS40UB>a+V#([B;Xe\\]
;+LVR3Zde=X3fGPQ(X>dJ)9R8$
`endprotected
endmodule



